magic
tech sky130A
magscale 1 2
timestamp 1745257087
<< checkpaint >>
rect -3932 -3108 10832 14396
<< viali >>
rect 1593 9061 1627 9095
rect 5365 9061 5399 9095
rect 4353 8993 4387 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 4445 8925 4479 8959
rect 5181 8925 5215 8959
rect 1869 8789 1903 8823
rect 4813 8789 4847 8823
rect 5365 8585 5399 8619
rect 4721 8449 4755 8483
rect 5181 8449 5215 8483
rect 4905 8381 4939 8415
rect 4537 8313 4571 8347
rect 1409 7837 1443 7871
rect 5181 7837 5215 7871
rect 1593 7701 1627 7735
rect 5365 7701 5399 7735
rect 4169 7497 4203 7531
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 3801 7361 3835 7395
rect 2973 7293 3007 7327
rect 3893 7293 3927 7327
rect 2973 7157 3007 7191
rect 3341 7157 3375 7191
rect 4077 6817 4111 6851
rect 4353 6817 4387 6851
rect 1409 6749 1443 6783
rect 3985 6749 4019 6783
rect 5181 6749 5215 6783
rect 1593 6613 1627 6647
rect 5365 6613 5399 6647
rect 2237 6409 2271 6443
rect 2053 6273 2087 6307
rect 4169 6273 4203 6307
rect 3617 6205 3651 6239
rect 4077 6205 4111 6239
rect 3709 6137 3743 6171
rect 4353 6069 4387 6103
rect 2053 5865 2087 5899
rect 1685 5797 1719 5831
rect 3525 5797 3559 5831
rect 1777 5729 1811 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 3341 5661 3375 5695
rect 3801 5321 3835 5355
rect 4077 5253 4111 5287
rect 1409 5185 1443 5219
rect 1593 5185 1627 5219
rect 1685 5185 1719 5219
rect 2329 5185 2363 5219
rect 2513 5185 2547 5219
rect 3709 5185 3743 5219
rect 3893 5185 3927 5219
rect 4261 5185 4295 5219
rect 5181 5185 5215 5219
rect 2421 5117 2455 5151
rect 4445 5117 4479 5151
rect 1593 5049 1627 5083
rect 1869 4981 1903 5015
rect 5365 4981 5399 5015
rect 3157 4777 3191 4811
rect 3801 4777 3835 4811
rect 4261 4777 4295 4811
rect 2789 4641 2823 4675
rect 3893 4641 3927 4675
rect 2973 4573 3007 4607
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 1409 4097 1443 4131
rect 5181 4097 5215 4131
rect 1593 3961 1627 3995
rect 5365 3893 5399 3927
rect 3433 3689 3467 3723
rect 3341 3621 3375 3655
rect 3203 3553 3237 3587
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 2881 3145 2915 3179
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 1593 2601 1627 2635
rect 1869 2533 1903 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2958 9092 2964 9104
rect 1627 9064 2964 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 3108 8996 4353 9024
rect 3108 8984 3114 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 1688 8888 1716 8919
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 3752 8928 4445 8956
rect 3752 8916 3758 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4764 8928 5181 8956
rect 4764 8916 4770 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 900 8860 1716 8888
rect 900 8848 906 8860
rect 1854 8780 1860 8832
rect 1912 8780 1918 8832
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 5166 8820 5172 8832
rect 4847 8792 5172 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5442 8616 5448 8628
rect 5399 8588 5448 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 4396 8452 4721 8480
rect 4396 8440 4402 8452
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4856 8452 5181 8480
rect 4856 8440 4862 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4304 8384 4905 8412
rect 4304 8372 4310 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 4522 8304 4528 8356
rect 4580 8304 4586 8356
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1670 7732 1676 7744
rect 1627 7704 1676 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 4154 7488 4160 7540
rect 4212 7488 4218 7540
rect 1854 7420 1860 7472
rect 1912 7460 1918 7472
rect 1912 7432 3188 7460
rect 1912 7420 1918 7432
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3160 7401 3188 7432
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 1728 7296 2973 7324
rect 1728 7284 1734 7296
rect 2961 7293 2973 7296
rect 3007 7324 3019 7327
rect 3804 7324 3832 7355
rect 3007 7296 3832 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3878 7284 3884 7336
rect 3936 7284 3942 7336
rect 2958 7148 2964 7200
rect 3016 7148 3022 7200
rect 3326 7148 3332 7200
rect 3384 7148 3390 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4246 6848 4252 6860
rect 4111 6820 4252 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 5074 6848 5080 6860
rect 4387 6820 5080 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4212 6752 5181 6780
rect 4212 6740 4218 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 1578 6604 1584 6656
rect 1636 6644 1642 6656
rect 2866 6644 2872 6656
rect 1636 6616 2872 6644
rect 1636 6604 1642 6616
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 4154 6440 4160 6452
rect 2271 6412 4160 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4522 6304 4528 6316
rect 4203 6276 4528 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 2056 6236 2084 6267
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 2056 6208 3617 6236
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3697 6171 3755 6177
rect 3697 6168 3709 6171
rect 3384 6140 3709 6168
rect 3384 6128 3390 6140
rect 3697 6137 3709 6140
rect 3743 6137 3755 6171
rect 3697 6131 3755 6137
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 4614 6100 4620 6112
rect 4387 6072 4620 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 4062 5896 4068 5908
rect 2087 5868 4068 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 1670 5788 1676 5840
rect 1728 5788 1734 5840
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 4798 5828 4804 5840
rect 3559 5800 4804 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 1811 5732 3004 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2976 5704 3004 5732
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 1854 5652 1860 5704
rect 1912 5652 1918 5704
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 3016 5664 3341 5692
rect 3016 5652 3022 5664
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3786 5556 3792 5568
rect 3384 5528 3792 5556
rect 3384 5516 3390 5528
rect 3786 5516 3792 5528
rect 3844 5556 3850 5568
rect 4062 5556 4068 5568
rect 3844 5528 4068 5556
rect 3844 5516 3850 5528
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 3050 5352 3056 5364
rect 1412 5324 3056 5352
rect 1412 5225 1440 5324
rect 3050 5312 3056 5324
rect 3108 5352 3114 5364
rect 3234 5352 3240 5364
rect 3108 5324 3240 5352
rect 3108 5312 3114 5324
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 4706 5352 4712 5364
rect 3835 5324 4712 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 4065 5287 4123 5293
rect 4065 5284 4077 5287
rect 1596 5256 4077 5284
rect 1596 5225 1624 5256
rect 4065 5253 4077 5256
rect 4111 5253 4123 5287
rect 4065 5247 4123 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1688 5148 1716 5179
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 2314 5216 2320 5228
rect 1912 5188 2320 5216
rect 1912 5176 1918 5188
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2958 5216 2964 5228
rect 2547 5188 2964 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3697 5219 3755 5225
rect 3697 5216 3709 5219
rect 3200 5188 3709 5216
rect 3200 5176 3206 5188
rect 3697 5185 3709 5188
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4212 5188 4261 5216
rect 4212 5176 4218 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 900 5120 1716 5148
rect 2409 5151 2467 5157
rect 900 5108 906 5120
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 3896 5148 3924 5176
rect 2455 5120 3924 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 4120 5120 4445 5148
rect 4120 5108 4126 5120
rect 4433 5117 4445 5120
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 5184 5080 5212 5179
rect 1627 5052 5212 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 1857 5015 1915 5021
rect 1857 4981 1869 5015
rect 1903 5012 1915 5015
rect 3050 5012 3056 5024
rect 1903 4984 3056 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 3050 4972 3056 4984
rect 3108 5012 3114 5024
rect 4062 5012 4068 5024
rect 3108 4984 4068 5012
rect 3108 4972 3114 4984
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 4246 4768 4252 4820
rect 4304 4768 4310 4820
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2777 4675 2835 4681
rect 2777 4672 2789 4675
rect 2372 4644 2789 4672
rect 2372 4632 2378 4644
rect 2777 4641 2789 4644
rect 2823 4641 2835 4675
rect 2777 4635 2835 4641
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3568 4644 3893 4672
rect 3568 4632 3574 4644
rect 3881 4641 3893 4644
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 2958 4564 2964 4616
rect 3016 4564 3022 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 3694 3992 3700 4004
rect 1627 3964 3700 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 4338 3720 4344 3732
rect 3467 3692 4344 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 3016 3624 3341 3652
rect 3016 3612 3022 3624
rect 3329 3621 3341 3624
rect 3375 3652 3387 3655
rect 3786 3652 3792 3664
rect 3375 3624 3792 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 3191 3587 3249 3593
rect 3191 3553 3203 3587
rect 3237 3584 3249 3587
rect 3694 3584 3700 3596
rect 3237 3556 3700 3584
rect 3237 3553 3249 3556
rect 3191 3547 3249 3553
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 3510 3476 3516 3528
rect 3568 3476 3574 3528
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3234 3176 3240 3188
rect 2915 3148 3240 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3050 3108 3056 3120
rect 2792 3080 3056 3108
rect 2792 3049 2820 3080
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3510 2632 3516 2644
rect 1627 2604 3516 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 3970 2564 3976 2576
rect 1903 2536 3976 2564
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 2964 9052 3016 9104
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 3056 8984 3108 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 848 8848 900 8900
rect 3700 8916 3752 8968
rect 4712 8916 4764 8968
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 5172 8780 5224 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 5448 8576 5500 8628
rect 4344 8440 4396 8492
rect 4804 8440 4856 8492
rect 4252 8372 4304 8424
rect 4528 8347 4580 8356
rect 4528 8313 4537 8347
rect 4537 8313 4571 8347
rect 4571 8313 4580 8347
rect 4528 8304 4580 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 848 7828 900 7880
rect 4160 7828 4212 7880
rect 1676 7692 1728 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 1860 7420 1912 7472
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 1676 7284 1728 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 4252 6808 4304 6860
rect 5080 6808 5132 6860
rect 848 6740 900 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4160 6740 4212 6792
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2872 6604 2924 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 4160 6400 4212 6452
rect 4528 6264 4580 6316
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 3332 6128 3384 6180
rect 4620 6060 4672 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 4068 5856 4120 5908
rect 1676 5831 1728 5840
rect 1676 5797 1685 5831
rect 1685 5797 1719 5831
rect 1719 5797 1728 5831
rect 1676 5788 1728 5797
rect 4804 5788 4856 5840
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2964 5652 3016 5704
rect 3332 5516 3384 5568
rect 3792 5516 3844 5568
rect 4068 5516 4120 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 3056 5312 3108 5364
rect 3240 5312 3292 5364
rect 4712 5312 4764 5364
rect 848 5108 900 5160
rect 1860 5176 1912 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 2964 5176 3016 5228
rect 3148 5176 3200 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4160 5176 4212 5228
rect 4068 5108 4120 5160
rect 3056 4972 3108 5024
rect 4068 4972 4120 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3700 4768 3752 4820
rect 4252 4811 4304 4820
rect 4252 4777 4261 4811
rect 4261 4777 4295 4811
rect 4295 4777 4304 4811
rect 4252 4768 4304 4777
rect 2320 4632 2372 4684
rect 3516 4632 3568 4684
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 848 4088 900 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 3700 3952 3752 4004
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 4344 3680 4396 3732
rect 2964 3612 3016 3664
rect 3792 3612 3844 3664
rect 3700 3544 3752 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 3240 3136 3292 3188
rect 3056 3068 3108 3120
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 3516 2592 3568 2644
rect 3976 2524 4028 2576
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 5446 10432 5502 10441
rect 5446 10367 5502 10376
rect 1412 8974 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 2964 9104 3016 9110
rect 5356 9104 5408 9110
rect 2964 9046 3016 9052
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 1400 8968 1452 8974
rect 846 8936 902 8945
rect 1400 8910 1452 8916
rect 846 8871 848 8880
rect 900 8871 902 8880
rect 848 8842 900 8848
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 900 7848 902 7857
rect 846 7783 902 7792
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7342 1716 7686
rect 1872 7478 1900 8774
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1596 5710 1624 6598
rect 1688 5846 1716 7278
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1872 5710 1900 7414
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2884 6662 2912 7346
rect 2976 7206 3004 9046
rect 3056 9036 3108 9042
rect 5354 9007 5410 9016
rect 3056 8978 3108 8984
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2976 5710 3004 7142
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 1872 5234 1900 5646
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2976 5234 3004 5646
rect 3068 5370 3096 8978
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6186 3372 7142
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3344 5574 3372 6122
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 848 5160 900 5166
rect 846 5128 848 5137
rect 900 5128 902 5137
rect 846 5063 902 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2332 4690 2360 5170
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2976 4622 3004 5170
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 846 3768 902 3777
rect 1950 3771 2258 3780
rect 846 3703 902 3712
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2976 3058 3004 3606
rect 3068 3534 3096 4966
rect 3160 4826 3188 5170
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 3126 3096 3470
rect 3252 3194 3280 5306
rect 3712 4826 3740 8910
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 3534 3556 4626
rect 3712 4010 3740 4762
rect 3804 4622 3832 5510
rect 3896 5234 3924 7278
rect 4264 6866 4292 8366
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3712 3602 3740 3946
rect 3804 3670 3832 4558
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3528 2650 3556 3470
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3988 2582 4016 6734
rect 4172 6458 4200 6734
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5914 4108 6190
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5250 4108 5510
rect 4080 5234 4200 5250
rect 4080 5228 4212 5234
rect 4080 5222 4160 5228
rect 4160 5170 4212 5176
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 5030 4108 5102
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4622 4108 4966
rect 4264 4826 4292 6802
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4356 3738 4384 8434
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4540 6322 4568 8298
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4632 2446 4660 6054
rect 4724 5370 4752 8910
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4816 5846 4844 8434
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 5092 2446 5120 6802
rect 5184 4146 5212 8774
rect 5460 8634 5488 10367
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6361 5396 6598
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 5446 10376 5502 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 846 8900 902 8936
rect 846 8880 848 8900
rect 848 8880 900 8900
rect 900 8880 902 8900
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 846 6432 902 6488
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 5354 9016 5410 9052
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 846 5108 848 5128
rect 848 5108 900 5128
rect 900 5108 902 5128
rect 846 5072 902 5108
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 846 3712 902 3768
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 5441 10434 5507 10437
rect 6100 10434 6900 10464
rect 5441 10432 6900 10434
rect 5441 10376 5446 10432
rect 5502 10376 6900 10432
rect 5441 10374 6900 10376
rect 5441 10371 5507 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_
timestamp 0
transform -1 0 2116 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _13_
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 0
transform -1 0 4140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 0
transform -1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 0
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _17_
timestamp 0
transform -1 0 4508 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 0
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 0
transform 1 0 4232 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _20_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _21_
timestamp 0
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform -1 0 4968 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform -1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 0
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 0
transform -1 0 3588 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_33
timestamp 0
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_45
timestamp 0
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_30
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_42
timestamp 0
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 0
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_35
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_9
timestamp 0
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_16
timestamp 0
transform 1 0 2576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_37
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_11
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_23
timestamp 0
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_9
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_13
timestamp 0
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_25
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_36
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 0
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_36
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_26
timestamp 0
transform 1 0 3496 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_34
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_46
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_35
timestamp 0
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_42
timestamp 0
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 0
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 3174 5134 3174 5134 4 _00_
rlabel metal1 s 3082 5882 3082 5882 4 _01_
rlabel metal1 s 3542 6154 3542 6154 4 _02_
rlabel metal1 s 2070 6256 2070 6256 4 _03_
rlabel metal1 s 1426 5270 1426 5270 4 _04_
rlabel metal1 s 1610 5236 1610 5236 4 _05_
rlabel metal1 s 4186 6834 4186 6834 4 _06_
rlabel metal1 s 3910 3706 3910 3706 4 _07_
rlabel metal1 s 4370 6290 4370 6290 4 _08_
rlabel metal2 s 3174 4998 3174 4998 4 _09_
rlabel metal3 s 1050 10404 1050 10404 4 in[0]
rlabel metal3 s 0 8984 800 9104 4 in[1]
port 4 nsew
rlabel metal3 s 0 7624 800 7744 4 in[2]
port 5 nsew
rlabel metal3 s 0 6264 800 6384 4 in[3]
port 6 nsew
rlabel metal3 s 0 4904 800 5024 4 in[4]
port 7 nsew
rlabel metal3 s 0 3544 800 3664 4 in[5]
port 8 nsew
rlabel metal3 s 0 2184 800 2304 4 in[6]
port 9 nsew
rlabel metal3 s 1188 884 1188 884 4 in[7]
rlabel metal1 s 3174 5678 3174 5678 4 net1
rlabel metal1 s 4278 5338 4278 5338 4 net10
rlabel metal2 s 4186 7684 4186 7684 4 net11
rlabel metal1 s 3220 6426 3220 6426 4 net12
rlabel metal1 s 5198 5134 5198 5134 4 net13
rlabel metal1 s 5014 8806 5014 8806 4 net14
rlabel metal2 s 4646 4250 4646 4250 4 net15
rlabel metal1 s 4738 6834 4738 6834 4 net16
rlabel metal1 s 2116 5202 2116 5202 4 net2
rlabel metal1 s 1656 7718 1656 7718 4 net3
rlabel metal1 s 2254 6630 2254 6630 4 net4
rlabel metal1 s 4278 5134 4278 5134 4 net5
rlabel metal1 s 3772 4794 3772 4794 4 net6
rlabel metal2 s 3542 3060 3542 3060 4 net7
rlabel metal1 s 2944 2550 2944 2550 4 net8
rlabel metal1 s 4186 5814 4186 5814 4 net9
rlabel metal1 s 5428 8602 5428 8602 4 out[0]
rlabel metal3 s 5382 9061 5382 9061 4 out[1]
rlabel metal3 s 5382 7701 5382 7701 4 out[2]
rlabel metal2 s 5382 6477 5382 6477 4 out[3]
rlabel metal3 s 5382 4981 5382 4981 4 out[4]
rlabel metal2 s 5382 3757 5382 3757 4 out[5]
rlabel metal3 s 4830 2261 4830 2261 4 out[6]
rlabel metal2 s 5474 1615 5474 1615 4 out[7]
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 10344 800 10464 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 400 9044 400 9044 0 FreeSans 600 0 0 0 in[1]
flabel metal3 s 400 7684 400 7684 0 FreeSans 600 0 0 0 in[2]
flabel metal3 s 400 6324 400 6324 0 FreeSans 600 0 0 0 in[3]
flabel metal3 s 400 4964 400 4964 0 FreeSans 600 0 0 0 in[4]
flabel metal3 s 400 3604 400 3604 0 FreeSans 600 0 0 0 in[5]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 0 824 800 944 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 600 0 0 0 out[2]
port 13 nsew
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 6100 824 6900 944 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
