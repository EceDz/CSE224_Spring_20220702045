magic
tech sky130A
magscale 1 2
timestamp 1747316550
<< viali >>
rect 5365 17289 5399 17323
rect 15301 17289 15335 17323
rect 18521 17289 18555 17323
rect 4629 17221 4663 17255
rect 8493 17221 8527 17255
rect 11989 17221 12023 17255
rect 15669 17221 15703 17255
rect 15945 17221 15979 17255
rect 15439 17187 15473 17221
rect 4445 17153 4479 17187
rect 7481 17153 7515 17187
rect 7665 17153 7699 17187
rect 7757 17153 7791 17187
rect 7849 17153 7883 17187
rect 13737 17153 13771 17187
rect 14749 17153 14783 17187
rect 7297 17085 7331 17119
rect 11713 17085 11747 17119
rect 15025 17085 15059 17119
rect 4997 17017 5031 17051
rect 8125 17017 8159 17051
rect 2881 16949 2915 16983
rect 4261 16949 4295 16983
rect 14381 16949 14415 16983
rect 14657 16949 14691 16983
rect 15485 16949 15519 16983
rect 2605 16745 2639 16779
rect 2237 16609 2271 16643
rect 2973 16609 3007 16643
rect 4721 16609 4755 16643
rect 6929 16609 6963 16643
rect 12357 16609 12391 16643
rect 14197 16609 14231 16643
rect 2329 16541 2363 16575
rect 3157 16541 3191 16575
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 5641 16541 5675 16575
rect 5825 16541 5859 16575
rect 6009 16541 6043 16575
rect 7205 16541 7239 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 12909 16541 12943 16575
rect 13277 16541 13311 16575
rect 14381 16541 14415 16575
rect 5365 16473 5399 16507
rect 7113 16473 7147 16507
rect 12081 16473 12115 16507
rect 12541 16473 12575 16507
rect 13737 16473 13771 16507
rect 14565 16473 14599 16507
rect 15209 16473 15243 16507
rect 3249 16405 3283 16439
rect 4997 16405 5031 16439
rect 5917 16405 5951 16439
rect 6285 16405 6319 16439
rect 11897 16405 11931 16439
rect 13369 16405 13403 16439
rect 14933 16405 14967 16439
rect 18521 16405 18555 16439
rect 14841 16201 14875 16235
rect 15117 16201 15151 16235
rect 4169 16133 4203 16167
rect 5917 16133 5951 16167
rect 13277 16065 13311 16099
rect 15025 16065 15059 16099
rect 15301 16065 15335 16099
rect 6193 15997 6227 16031
rect 13001 15997 13035 16031
rect 15485 15929 15519 15963
rect 3065 15861 3099 15895
rect 11529 15861 11563 15895
rect 14013 15861 14047 15895
rect 14565 15861 14599 15895
rect 15393 15861 15427 15895
rect 15761 15861 15795 15895
rect 3617 15657 3651 15691
rect 7849 15657 7883 15691
rect 10057 15657 10091 15691
rect 11253 15657 11287 15691
rect 14105 15657 14139 15691
rect 7665 15589 7699 15623
rect 11529 15589 11563 15623
rect 1869 15521 1903 15555
rect 6285 15521 6319 15555
rect 7481 15521 7515 15555
rect 12173 15521 12207 15555
rect 1409 15453 1443 15487
rect 5273 15453 5307 15487
rect 5457 15453 5491 15487
rect 5733 15453 5767 15487
rect 5825 15453 5859 15487
rect 10609 15453 10643 15487
rect 10793 15453 10827 15487
rect 11437 15453 11471 15487
rect 11713 15453 11747 15487
rect 11805 15453 11839 15487
rect 14381 15453 14415 15487
rect 2145 15385 2179 15419
rect 3985 15385 4019 15419
rect 4537 15385 4571 15419
rect 4721 15385 4755 15419
rect 4905 15385 4939 15419
rect 5641 15385 5675 15419
rect 7205 15385 7239 15419
rect 7833 15385 7867 15419
rect 8033 15385 8067 15419
rect 10517 15385 10551 15419
rect 13829 15385 13863 15419
rect 14657 15385 14691 15419
rect 1593 15317 1627 15351
rect 4353 15317 4387 15351
rect 5089 15317 5123 15351
rect 5365 15317 5399 15351
rect 6653 15317 6687 15351
rect 10609 15317 10643 15351
rect 14289 15317 14323 15351
rect 14473 15317 14507 15351
rect 15301 15317 15335 15351
rect 18521 15317 18555 15351
rect 10793 15113 10827 15147
rect 13997 15113 14031 15147
rect 15209 15113 15243 15147
rect 15761 15113 15795 15147
rect 1593 15045 1627 15079
rect 5181 15045 5215 15079
rect 5825 15045 5859 15079
rect 9489 15045 9523 15079
rect 9689 15045 9723 15079
rect 14197 15045 14231 15079
rect 5641 14977 5675 15011
rect 5917 14977 5951 15011
rect 10057 14977 10091 15011
rect 10734 14977 10768 15011
rect 15025 14977 15059 15011
rect 15301 14977 15335 15011
rect 15853 14977 15887 15011
rect 6653 14909 6687 14943
rect 10517 14909 10551 14943
rect 11253 14909 11287 14943
rect 11713 14909 11747 14943
rect 15393 14909 15427 14943
rect 5641 14841 5675 14875
rect 2421 14773 2455 14807
rect 5549 14773 5583 14807
rect 9321 14773 9355 14807
rect 9505 14773 9539 14807
rect 10609 14773 10643 14807
rect 11161 14773 11195 14807
rect 13645 14773 13679 14807
rect 13829 14773 13863 14807
rect 14013 14773 14047 14807
rect 14657 14773 14691 14807
rect 15577 14773 15611 14807
rect 2237 14569 2271 14603
rect 4169 14569 4203 14603
rect 6653 14569 6687 14603
rect 9781 14569 9815 14603
rect 2605 14501 2639 14535
rect 12633 14501 12667 14535
rect 18337 14501 18371 14535
rect 3433 14433 3467 14467
rect 12357 14433 12391 14467
rect 15485 14433 15519 14467
rect 2145 14365 2179 14399
rect 2237 14365 2271 14399
rect 2697 14365 2731 14399
rect 2973 14365 3007 14399
rect 4905 14365 4939 14399
rect 8401 14365 8435 14399
rect 12541 14365 12575 14399
rect 12725 14365 12759 14399
rect 16037 14365 16071 14399
rect 18521 14365 18555 14399
rect 4537 14297 4571 14331
rect 8125 14297 8159 14331
rect 16313 14297 16347 14331
rect 1869 14229 1903 14263
rect 6009 14229 6043 14263
rect 17785 14229 17819 14263
rect 18245 14229 18279 14263
rect 4169 14025 4203 14059
rect 6577 14025 6611 14059
rect 6745 14025 6779 14059
rect 8401 14025 8435 14059
rect 11529 14025 11563 14059
rect 13369 14025 13403 14059
rect 15945 14025 15979 14059
rect 17417 14025 17451 14059
rect 18061 14025 18095 14059
rect 3893 13957 3927 13991
rect 5641 13957 5675 13991
rect 6377 13957 6411 13991
rect 8125 13957 8159 13991
rect 11681 13957 11715 13991
rect 11897 13957 11931 13991
rect 14105 13957 14139 13991
rect 3525 13889 3559 13923
rect 3801 13889 3835 13923
rect 3985 13889 4019 13923
rect 5917 13889 5951 13923
rect 7021 13889 7055 13923
rect 7205 13889 7239 13923
rect 7757 13889 7791 13923
rect 10241 13889 10275 13923
rect 10517 13889 10551 13923
rect 13093 13889 13127 13923
rect 13461 13889 13495 13923
rect 13829 13889 13863 13923
rect 15853 13889 15887 13923
rect 16129 13889 16163 13923
rect 17944 13889 17978 13923
rect 2605 13821 2639 13855
rect 6929 13821 6963 13855
rect 7297 13821 7331 13855
rect 10149 13821 10183 13855
rect 15577 13821 15611 13855
rect 15761 13821 15795 13855
rect 17141 13821 17175 13855
rect 18153 13821 18187 13855
rect 18429 13821 18463 13855
rect 6561 13685 6595 13719
rect 11713 13685 11747 13719
rect 12265 13685 12299 13719
rect 17785 13685 17819 13719
rect 8125 13481 8159 13515
rect 17693 13481 17727 13515
rect 18061 13481 18095 13515
rect 4721 13345 4755 13379
rect 6469 13345 6503 13379
rect 3893 13277 3927 13311
rect 4445 13277 4479 13311
rect 6745 13277 6779 13311
rect 6929 13277 6963 13311
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 8493 13277 8527 13311
rect 10241 13277 10275 13311
rect 10609 13277 10643 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13185 13277 13219 13311
rect 15301 13277 15335 13311
rect 6193 13209 6227 13243
rect 7849 13209 7883 13243
rect 10517 13209 10551 13243
rect 13461 13209 13495 13243
rect 15577 13209 15611 13243
rect 17325 13209 17359 13243
rect 4077 13141 4111 13175
rect 4629 13141 4663 13175
rect 6837 13141 6871 13175
rect 7389 13141 7423 13175
rect 18521 13141 18555 13175
rect 2789 12937 2823 12971
rect 18429 12937 18463 12971
rect 3709 12869 3743 12903
rect 6469 12869 6503 12903
rect 11129 12869 11163 12903
rect 11345 12869 11379 12903
rect 2881 12801 2915 12835
rect 3525 12801 3559 12835
rect 3617 12801 3651 12835
rect 7021 12801 7055 12835
rect 7573 12801 7607 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 10701 12801 10735 12835
rect 12265 12801 12299 12835
rect 13737 12801 13771 12835
rect 16681 12801 16715 12835
rect 7849 12733 7883 12767
rect 8125 12733 8159 12767
rect 10241 12733 10275 12767
rect 16221 12733 16255 12767
rect 16957 12733 16991 12767
rect 3065 12665 3099 12699
rect 7205 12665 7239 12699
rect 10701 12665 10735 12699
rect 13921 12665 13955 12699
rect 9597 12597 9631 12631
rect 10977 12597 11011 12631
rect 11161 12597 11195 12631
rect 11805 12597 11839 12631
rect 1961 12393 1995 12427
rect 2421 12393 2455 12427
rect 5549 12393 5583 12427
rect 10793 12393 10827 12427
rect 14473 12393 14507 12427
rect 14749 12393 14783 12427
rect 2605 12325 2639 12359
rect 5733 12257 5767 12291
rect 6285 12257 6319 12291
rect 16129 12257 16163 12291
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 5825 12189 5859 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 14657 12189 14691 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 16773 12189 16807 12223
rect 17141 12189 17175 12223
rect 17417 12189 17451 12223
rect 17693 12189 17727 12223
rect 2237 12121 2271 12155
rect 3801 12121 3835 12155
rect 8033 12121 8067 12155
rect 12725 12121 12759 12155
rect 2437 12053 2471 12087
rect 2973 12053 3007 12087
rect 4077 12053 4111 12087
rect 4353 12053 4387 12087
rect 4813 12053 4847 12087
rect 11897 12053 11931 12087
rect 12265 12053 12299 12087
rect 13093 12053 13127 12087
rect 13461 12053 13495 12087
rect 15209 12053 15243 12087
rect 15853 12053 15887 12087
rect 17049 12053 17083 12087
rect 17325 12053 17359 12087
rect 18521 12053 18555 12087
rect 8309 11849 8343 11883
rect 12265 11849 12299 11883
rect 14013 11849 14047 11883
rect 14657 11849 14691 11883
rect 14841 11849 14875 11883
rect 6837 11781 6871 11815
rect 16037 11781 16071 11815
rect 2605 11713 2639 11747
rect 4537 11713 4571 11747
rect 6561 11713 6595 11747
rect 8401 11713 8435 11747
rect 10425 11713 10459 11747
rect 11345 11713 11379 11747
rect 11933 11713 11967 11747
rect 12265 11713 12299 11747
rect 12449 11713 12483 11747
rect 12725 11713 12759 11747
rect 15577 11713 15611 11747
rect 16129 11713 16163 11747
rect 16497 11713 16531 11747
rect 8677 11645 8711 11679
rect 11529 11645 11563 11679
rect 11621 11645 11655 11679
rect 15209 11645 15243 11679
rect 15853 11645 15887 11679
rect 2789 11577 2823 11611
rect 10149 11577 10183 11611
rect 11253 11577 11287 11611
rect 15577 11577 15611 11611
rect 15669 11577 15703 11611
rect 3157 11509 3191 11543
rect 4721 11509 4755 11543
rect 10241 11509 10275 11543
rect 11069 11509 11103 11543
rect 12081 11509 12115 11543
rect 14841 11509 14875 11543
rect 6837 11305 6871 11339
rect 7113 11305 7147 11339
rect 10701 11305 10735 11339
rect 11345 11305 11379 11339
rect 11713 11305 11747 11339
rect 14933 11305 14967 11339
rect 17325 11305 17359 11339
rect 4905 11237 4939 11271
rect 6561 11237 6595 11271
rect 17141 11237 17175 11271
rect 9045 11169 9079 11203
rect 9505 11169 9539 11203
rect 10885 11169 10919 11203
rect 11897 11169 11931 11203
rect 13921 11169 13955 11203
rect 15853 11169 15887 11203
rect 4721 11101 4755 11135
rect 6377 11101 6411 11135
rect 6653 11101 6687 11135
rect 7205 11101 7239 11135
rect 8769 11101 8803 11135
rect 9137 11101 9171 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 10701 11101 10735 11135
rect 10977 11101 11011 11135
rect 14105 11101 14139 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 17049 11101 17083 11135
rect 10425 11033 10459 11067
rect 12173 11033 12207 11067
rect 14197 11033 14231 11067
rect 14565 11033 14599 11067
rect 15669 11033 15703 11067
rect 17309 11033 17343 11067
rect 17509 11033 17543 11067
rect 18521 11033 18555 11067
rect 16221 10965 16255 10999
rect 9045 10761 9079 10795
rect 10793 10761 10827 10795
rect 11345 10761 11379 10795
rect 11897 10761 11931 10795
rect 11529 10693 11563 10727
rect 11713 10693 11747 10727
rect 12449 10693 12483 10727
rect 16957 10693 16991 10727
rect 2697 10625 2731 10659
rect 6377 10625 6411 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 8769 10625 8803 10659
rect 9045 10625 9079 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 17141 10625 17175 10659
rect 2973 10557 3007 10591
rect 12081 10557 12115 10591
rect 7665 10489 7699 10523
rect 8953 10489 8987 10523
rect 4445 10421 4479 10455
rect 6561 10421 6595 10455
rect 7941 10421 7975 10455
rect 9321 10421 9355 10455
rect 13921 10421 13955 10455
rect 17233 10421 17267 10455
rect 10977 10081 11011 10115
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 18521 10013 18555 10047
rect 6101 9945 6135 9979
rect 6469 9945 6503 9979
rect 8677 9945 8711 9979
rect 9229 9945 9263 9979
rect 5733 9877 5767 9911
rect 12909 9673 12943 9707
rect 4997 9605 5031 9639
rect 9413 9605 9447 9639
rect 7113 9537 7147 9571
rect 7389 9537 7423 9571
rect 7665 9537 7699 9571
rect 10057 9537 10091 9571
rect 12357 9537 12391 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 2973 9469 3007 9503
rect 3249 9469 3283 9503
rect 7205 9469 7239 9503
rect 9689 9469 9723 9503
rect 7297 9401 7331 9435
rect 12357 9401 12391 9435
rect 6837 9333 6871 9367
rect 7573 9333 7607 9367
rect 11989 9333 12023 9367
rect 6285 9129 6319 9163
rect 6745 9129 6779 9163
rect 9781 9129 9815 9163
rect 10885 9129 10919 9163
rect 10977 9129 11011 9163
rect 13737 9129 13771 9163
rect 18061 9129 18095 9163
rect 8217 9061 8251 9095
rect 9045 9061 9079 9095
rect 11529 9061 11563 9095
rect 17049 9061 17083 9095
rect 9689 8993 9723 9027
rect 9940 8993 9974 9027
rect 10057 8993 10091 9027
rect 10425 8993 10459 9027
rect 11989 8993 12023 9027
rect 2605 8925 2639 8959
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 6837 8925 6871 8959
rect 7573 8925 7607 8959
rect 7757 8925 7791 8959
rect 8309 8925 8343 8959
rect 10977 8925 11011 8959
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 17417 8925 17451 8959
rect 18245 8925 18279 8959
rect 2697 8857 2731 8891
rect 3249 8857 3283 8891
rect 3985 8857 4019 8891
rect 7481 8857 7515 8891
rect 10517 8857 10551 8891
rect 10701 8857 10735 8891
rect 12265 8857 12299 8891
rect 17325 8857 17359 8891
rect 3065 8789 3099 8823
rect 3617 8789 3651 8823
rect 7665 8789 7699 8823
rect 8677 8789 8711 8823
rect 10149 8789 10183 8823
rect 14289 8789 14323 8823
rect 18429 8789 18463 8823
rect 3433 8585 3467 8619
rect 10609 8585 10643 8619
rect 11345 8585 11379 8619
rect 12541 8585 12575 8619
rect 13369 8585 13403 8619
rect 14197 8585 14231 8619
rect 4905 8517 4939 8551
rect 6377 8517 6411 8551
rect 8033 8517 8067 8551
rect 10057 8517 10091 8551
rect 12173 8517 12207 8551
rect 12357 8517 12391 8551
rect 18153 8517 18187 8551
rect 3617 8449 3651 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 9956 8439 9990 8473
rect 10251 8449 10285 8483
rect 12449 8449 12483 8483
rect 13001 8449 13035 8483
rect 13645 8449 13679 8483
rect 14105 8449 14139 8483
rect 14289 8449 14323 8483
rect 17417 8449 17451 8483
rect 1685 8381 1719 8415
rect 1961 8381 1995 8415
rect 4629 8381 4663 8415
rect 9781 8381 9815 8415
rect 11805 8381 11839 8415
rect 14565 8381 14599 8415
rect 4261 8313 4295 8347
rect 8401 8313 8435 8347
rect 9413 8313 9447 8347
rect 10241 8313 10275 8347
rect 10885 8313 10919 8347
rect 12725 8313 12759 8347
rect 12909 8313 12943 8347
rect 17509 8313 17543 8347
rect 18429 8245 18463 8279
rect 2145 8041 2179 8075
rect 2789 8041 2823 8075
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 13369 8041 13403 8075
rect 13553 8041 13587 8075
rect 17693 8041 17727 8075
rect 4261 7973 4295 8007
rect 6837 7973 6871 8007
rect 10333 7905 10367 7939
rect 12541 7905 12575 7939
rect 17969 7905 18003 7939
rect 3525 7837 3559 7871
rect 3801 7837 3835 7871
rect 4813 7837 4847 7871
rect 7113 7837 7147 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 17877 7837 17911 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 2605 7769 2639 7803
rect 2821 7769 2855 7803
rect 5089 7769 5123 7803
rect 6837 7769 6871 7803
rect 12265 7769 12299 7803
rect 14289 7769 14323 7803
rect 14933 7769 14967 7803
rect 2513 7701 2547 7735
rect 2973 7701 3007 7735
rect 4721 7701 4755 7735
rect 6561 7701 6595 7735
rect 7021 7701 7055 7735
rect 7389 7701 7423 7735
rect 10793 7701 10827 7735
rect 12909 7701 12943 7735
rect 13921 7701 13955 7735
rect 17325 7701 17359 7735
rect 18429 7701 18463 7735
rect 7849 7497 7883 7531
rect 10333 7497 10367 7531
rect 11069 7497 11103 7531
rect 12817 7497 12851 7531
rect 14933 7497 14967 7531
rect 17601 7497 17635 7531
rect 2697 7429 2731 7463
rect 10977 7429 11011 7463
rect 11529 7429 11563 7463
rect 17141 7429 17175 7463
rect 7941 7361 7975 7395
rect 8217 7361 8251 7395
rect 10425 7361 10459 7395
rect 10609 7361 10643 7395
rect 13553 7361 13587 7395
rect 16405 7361 16439 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 2421 7293 2455 7327
rect 4169 7293 4203 7327
rect 4445 7293 4479 7327
rect 4721 7293 4755 7327
rect 6193 7293 6227 7327
rect 10517 7293 10551 7327
rect 14289 7225 14323 7259
rect 14657 7225 14691 7259
rect 17417 7225 17451 7259
rect 17969 7225 18003 7259
rect 16773 7157 16807 7191
rect 17601 7157 17635 7191
rect 3525 6953 3559 6987
rect 8677 6953 8711 6987
rect 9505 6953 9539 6987
rect 11621 6953 11655 6987
rect 12449 6953 12483 6987
rect 12633 6953 12667 6987
rect 17141 6953 17175 6987
rect 17969 6953 18003 6987
rect 13553 6885 13587 6919
rect 3985 6817 4019 6851
rect 6561 6817 6595 6851
rect 9413 6817 9447 6851
rect 10057 6817 10091 6851
rect 11253 6817 11287 6851
rect 11437 6817 11471 6851
rect 13829 6817 13863 6851
rect 14565 6817 14599 6851
rect 15577 6817 15611 6851
rect 6009 6749 6043 6783
rect 6653 6749 6687 6783
rect 6929 6749 6963 6783
rect 7113 6749 7147 6783
rect 7389 6749 7423 6783
rect 9781 6749 9815 6783
rect 11337 6749 11371 6783
rect 11621 6749 11655 6783
rect 11769 6749 11803 6783
rect 11897 6749 11931 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 14289 6749 14323 6783
rect 14933 6749 14967 6783
rect 15025 6749 15059 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 18245 6749 18279 6783
rect 4261 6681 4295 6715
rect 6377 6681 6411 6715
rect 9505 6681 9539 6715
rect 12265 6681 12299 6715
rect 14749 6681 14783 6715
rect 15393 6681 15427 6715
rect 17417 6681 17451 6715
rect 3065 6613 3099 6647
rect 7021 6613 7055 6647
rect 7205 6613 7239 6647
rect 9689 6613 9723 6647
rect 10885 6613 10919 6647
rect 12449 6613 12483 6647
rect 12817 6613 12851 6647
rect 15945 6613 15979 6647
rect 18429 6613 18463 6647
rect 3801 6409 3835 6443
rect 3893 6409 3927 6443
rect 5917 6409 5951 6443
rect 9873 6409 9907 6443
rect 11913 6409 11947 6443
rect 12725 6409 12759 6443
rect 15301 6409 15335 6443
rect 17325 6409 17359 6443
rect 11713 6341 11747 6375
rect 13185 6341 13219 6375
rect 13829 6341 13863 6375
rect 15485 6341 15519 6375
rect 17141 6341 17175 6375
rect 4077 6273 4111 6307
rect 4169 6273 4203 6307
rect 4261 6273 4295 6307
rect 4537 6273 4571 6307
rect 4721 6273 4755 6307
rect 5733 6273 5767 6307
rect 9781 6273 9815 6307
rect 10241 6273 10275 6307
rect 13553 6273 13587 6307
rect 15393 6273 15427 6307
rect 15669 6273 15703 6307
rect 16037 6273 16071 6307
rect 16865 6273 16899 6307
rect 16957 6273 16991 6307
rect 17233 6273 17267 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 18153 6273 18187 6307
rect 18337 6273 18371 6307
rect 4905 6205 4939 6239
rect 17417 6205 17451 6239
rect 4445 6137 4479 6171
rect 5549 6137 5583 6171
rect 12357 6137 12391 6171
rect 15853 6137 15887 6171
rect 16865 6137 16899 6171
rect 18153 6137 18187 6171
rect 5181 6069 5215 6103
rect 11345 6069 11379 6103
rect 11897 6069 11931 6103
rect 12081 6069 12115 6103
rect 16129 6069 16163 6103
rect 2789 5865 2823 5899
rect 3525 5865 3559 5899
rect 4537 5865 4571 5899
rect 5825 5865 5859 5899
rect 8033 5865 8067 5899
rect 10793 5865 10827 5899
rect 11253 5865 11287 5899
rect 12817 5865 12851 5899
rect 13093 5865 13127 5899
rect 13277 5865 13311 5899
rect 15209 5865 15243 5899
rect 15577 5865 15611 5899
rect 17417 5865 17451 5899
rect 17877 5865 17911 5899
rect 5089 5797 5123 5831
rect 16313 5797 16347 5831
rect 2145 5729 2179 5763
rect 3157 5729 3191 5763
rect 14933 5729 14967 5763
rect 2329 5661 2363 5695
rect 2605 5661 2639 5695
rect 2789 5661 2823 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5457 5661 5491 5695
rect 13553 5661 13587 5695
rect 13921 5661 13955 5695
rect 16681 5661 16715 5695
rect 18245 5661 18279 5695
rect 4905 5593 4939 5627
rect 9965 5593 9999 5627
rect 10609 5593 10643 5627
rect 10809 5593 10843 5627
rect 13261 5593 13295 5627
rect 13461 5593 13495 5627
rect 13737 5593 13771 5627
rect 17049 5593 17083 5627
rect 2513 5525 2547 5559
rect 4445 5525 4479 5559
rect 10977 5525 11011 5559
rect 18429 5525 18463 5559
rect 2697 5321 2731 5355
rect 7481 5321 7515 5355
rect 10333 5321 10367 5355
rect 13645 5321 13679 5355
rect 13921 5321 13955 5355
rect 15853 5321 15887 5355
rect 16681 5321 16715 5355
rect 17049 5321 17083 5355
rect 17233 5321 17267 5355
rect 18153 5321 18187 5355
rect 2421 5253 2455 5287
rect 7297 5253 7331 5287
rect 8309 5253 8343 5287
rect 10149 5253 10183 5287
rect 10701 5253 10735 5287
rect 2605 5185 2639 5219
rect 3065 5185 3099 5219
rect 7389 5185 7423 5219
rect 7665 5185 7699 5219
rect 8033 5185 8067 5219
rect 10057 5185 10091 5219
rect 10425 5185 10459 5219
rect 17785 5185 17819 5219
rect 16865 5117 16899 5151
rect 16957 5117 16991 5151
rect 17325 5117 17359 5151
rect 10149 5049 10183 5083
rect 2329 4981 2363 5015
rect 7849 4981 7883 5015
rect 13277 4981 13311 5015
rect 16129 4981 16163 5015
rect 3985 4777 4019 4811
rect 4353 4777 4387 4811
rect 7021 4777 7055 4811
rect 7205 4777 7239 4811
rect 8125 4777 8159 4811
rect 12541 4777 12575 4811
rect 16129 4777 16163 4811
rect 16589 4777 16623 4811
rect 17049 4777 17083 4811
rect 17233 4777 17267 4811
rect 10241 4709 10275 4743
rect 10793 4709 10827 4743
rect 12173 4709 12207 4743
rect 14657 4709 14691 4743
rect 15577 4709 15611 4743
rect 18153 4709 18187 4743
rect 6929 4641 6963 4675
rect 3801 4573 3835 4607
rect 6745 4573 6779 4607
rect 7021 4573 7055 4607
rect 7481 4573 7515 4607
rect 9965 4573 9999 4607
rect 10241 4573 10275 4607
rect 10609 4573 10643 4607
rect 12725 4573 12759 4607
rect 12909 4573 12943 4607
rect 13185 4573 13219 4607
rect 17417 4573 17451 4607
rect 18245 4573 18279 4607
rect 8769 4505 8803 4539
rect 8953 4505 8987 4539
rect 9689 4505 9723 4539
rect 11161 4505 11195 4539
rect 14933 4505 14967 4539
rect 15117 4505 15151 4539
rect 15301 4505 15335 4539
rect 17785 4505 17819 4539
rect 18429 4437 18463 4471
rect 2053 4233 2087 4267
rect 7389 4233 7423 4267
rect 8401 4233 8435 4267
rect 8661 4233 8695 4267
rect 11897 4233 11931 4267
rect 12633 4233 12667 4267
rect 17509 4233 17543 4267
rect 18035 4233 18069 4267
rect 4261 4165 4295 4199
rect 8861 4165 8895 4199
rect 11529 4165 11563 4199
rect 11745 4165 11779 4199
rect 13369 4165 13403 4199
rect 18245 4165 18279 4199
rect 1869 4097 1903 4131
rect 2237 4097 2271 4131
rect 6009 4097 6043 4131
rect 6377 4097 6411 4131
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 18337 4097 18371 4131
rect 2421 4029 2455 4063
rect 3985 4029 4019 4063
rect 9321 4029 9355 4063
rect 9597 4029 9631 4063
rect 11345 4029 11379 4063
rect 13737 4029 13771 4063
rect 6561 3961 6595 3995
rect 8493 3961 8527 3995
rect 1777 3893 1811 3927
rect 2697 3893 2731 3927
rect 8677 3893 8711 3927
rect 11713 3893 11747 3927
rect 12173 3893 12207 3927
rect 17877 3893 17911 3927
rect 18061 3893 18095 3927
rect 18429 3893 18463 3927
rect 1961 3689 1995 3723
rect 2973 3689 3007 3723
rect 3249 3689 3283 3723
rect 9137 3689 9171 3723
rect 17601 3689 17635 3723
rect 11345 3621 11379 3655
rect 12357 3621 12391 3655
rect 6745 3553 6779 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 3157 3485 3191 3519
rect 8769 3485 8803 3519
rect 11621 3485 11655 3519
rect 11713 3485 11747 3519
rect 11805 3485 11839 3519
rect 11897 3485 11931 3519
rect 12173 3485 12207 3519
rect 17785 3485 17819 3519
rect 18245 3485 18279 3519
rect 7021 3417 7055 3451
rect 8953 3417 8987 3451
rect 9153 3417 9187 3451
rect 9321 3349 9355 3383
rect 12081 3349 12115 3383
rect 12633 3349 12667 3383
rect 13001 3349 13035 3383
rect 17877 3349 17911 3383
rect 18429 3349 18463 3383
rect 10333 3145 10367 3179
rect 11713 3145 11747 3179
rect 12541 3145 12575 3179
rect 13185 3145 13219 3179
rect 14565 3145 14599 3179
rect 15025 3145 15059 3179
rect 8861 3077 8895 3111
rect 10609 3077 10643 3111
rect 11529 3077 11563 3111
rect 10885 3009 10919 3043
rect 11805 3009 11839 3043
rect 11897 3009 11931 3043
rect 12817 3009 12851 3043
rect 11253 2873 11287 2907
rect 6101 2805 6135 2839
rect 12081 2805 12115 2839
rect 6009 2601 6043 2635
rect 6653 2601 6687 2635
rect 11253 2601 11287 2635
rect 14749 2601 14783 2635
rect 14933 2533 14967 2567
rect 9505 2465 9539 2499
rect 14381 2465 14415 2499
rect 15393 2465 15427 2499
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 15117 2397 15151 2431
rect 15209 2397 15243 2431
rect 15301 2397 15335 2431
rect 18245 2397 18279 2431
rect 9137 2329 9171 2363
rect 9781 2329 9815 2363
rect 5641 2261 5675 2295
rect 7021 2261 7055 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 15654 17592 15660 17604
rect 7340 17564 15660 17592
rect 7340 17552 7346 17564
rect 15654 17552 15660 17564
rect 15712 17552 15718 17604
rect 1104 17434 18860 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 18860 17434
rect 1104 17360 18860 17382
rect 5353 17323 5411 17329
rect 5353 17320 5365 17323
rect 4632 17292 5365 17320
rect 4632 17261 4660 17292
rect 5353 17289 5365 17292
rect 5399 17320 5411 17323
rect 9766 17320 9772 17332
rect 5399 17292 9772 17320
rect 5399 17289 5411 17292
rect 5353 17283 5411 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 10560 17292 15301 17320
rect 10560 17280 10566 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 18506 17280 18512 17332
rect 18564 17280 18570 17332
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17221 4675 17255
rect 8478 17252 8484 17264
rect 4617 17215 4675 17221
rect 7668 17224 8484 17252
rect 7668 17193 7696 17224
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 9732 17224 11989 17252
rect 9732 17212 9738 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 13446 17252 13452 17264
rect 13202 17224 13452 17252
rect 11977 17215 12035 17221
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 15427 17221 15485 17227
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 7469 17187 7527 17193
rect 4479 17156 5028 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 3418 17008 3424 17060
rect 3476 17048 3482 17060
rect 5000 17057 5028 17156
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7484 17116 7512 17147
rect 7742 17144 7748 17196
rect 7800 17144 7806 17196
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 10594 17184 10600 17196
rect 7883 17156 10600 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 13722 17144 13728 17196
rect 13780 17144 13786 17196
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14424 17156 14749 17184
rect 14424 17144 14430 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15427 17187 15439 17221
rect 15473 17187 15485 17221
rect 15654 17212 15660 17264
rect 15712 17252 15718 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15712 17224 15945 17252
rect 15712 17212 15718 17224
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 15427 17184 15485 17187
rect 14737 17147 14795 17153
rect 15028 17181 15485 17184
rect 15028 17156 15484 17181
rect 11606 17116 11612 17128
rect 7340 17088 7512 17116
rect 8036 17088 11612 17116
rect 7340 17076 7346 17088
rect 4985 17051 5043 17057
rect 3476 17020 4384 17048
rect 3476 17008 3482 17020
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16980 2927 16983
rect 3142 16980 3148 16992
rect 2915 16952 3148 16980
rect 2915 16949 2927 16952
rect 2869 16943 2927 16949
rect 3142 16940 3148 16952
rect 3200 16940 3206 16992
rect 4246 16940 4252 16992
rect 4304 16940 4310 16992
rect 4356 16980 4384 17020
rect 4985 17017 4997 17051
rect 5031 17048 5043 17051
rect 8036 17048 8064 17088
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 11698 17076 11704 17128
rect 11756 17076 11762 17128
rect 15028 17125 15056 17156
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 11808 17088 15025 17116
rect 5031 17020 8064 17048
rect 8113 17051 8171 17057
rect 5031 17017 5043 17020
rect 4985 17011 5043 17017
rect 8113 17017 8125 17051
rect 8159 17048 8171 17051
rect 10870 17048 10876 17060
rect 8159 17020 10876 17048
rect 8159 17017 8171 17020
rect 8113 17011 8171 17017
rect 10870 17008 10876 17020
rect 10928 17008 10934 17060
rect 11808 17048 11836 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 11624 17020 11836 17048
rect 11624 16980 11652 17020
rect 4356 16952 11652 16980
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 13262 16980 13268 16992
rect 11756 16952 13268 16980
rect 11756 16940 11762 16952
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 14642 16940 14648 16992
rect 14700 16940 14706 16992
rect 15473 16983 15531 16989
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 16758 16980 16764 16992
rect 15519 16952 16764 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 1104 16890 18860 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 18860 16890
rect 1104 16816 18860 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 1820 16748 2605 16776
rect 1820 16736 1826 16748
rect 2593 16745 2605 16748
rect 2639 16745 2651 16779
rect 2593 16739 2651 16745
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 13998 16776 14004 16788
rect 4304 16748 14004 16776
rect 4304 16736 4310 16748
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 3142 16708 3148 16720
rect 2240 16680 3148 16708
rect 2240 16649 2268 16680
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 3786 16668 3792 16720
rect 3844 16708 3850 16720
rect 3844 16680 6960 16708
rect 3844 16668 3850 16680
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16609 2283 16643
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2225 16603 2283 16609
rect 2332 16612 2973 16640
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2332 16581 2360 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 4709 16643 4767 16649
rect 4709 16609 4721 16643
rect 4755 16640 4767 16643
rect 5074 16640 5080 16652
rect 4755 16612 5080 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 2317 16575 2375 16581
rect 2317 16572 2329 16575
rect 1728 16544 2329 16572
rect 1728 16532 1734 16544
rect 2317 16541 2329 16544
rect 2363 16574 2375 16575
rect 3145 16575 3203 16581
rect 2363 16546 2397 16574
rect 2363 16541 2375 16546
rect 2317 16535 2375 16541
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3786 16572 3792 16584
rect 3191 16544 3792 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 5000 16581 5028 16612
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 6932 16649 6960 16680
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 14642 16708 14648 16720
rect 7524 16680 14648 16708
rect 7524 16668 7530 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 11698 16640 11704 16652
rect 6963 16612 11704 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16572 5043 16575
rect 5031 16544 5065 16572
rect 5031 16541 5043 16544
rect 4985 16535 5043 16541
rect 4338 16464 4344 16516
rect 4396 16504 4402 16516
rect 4816 16504 4844 16535
rect 5258 16532 5264 16584
rect 5316 16572 5322 16584
rect 7208 16581 7236 16612
rect 11698 16600 11704 16612
rect 11756 16640 11762 16652
rect 12345 16643 12403 16649
rect 11756 16612 12296 16640
rect 11756 16600 11762 16612
rect 5629 16575 5687 16581
rect 5629 16572 5641 16575
rect 5316 16544 5641 16572
rect 5316 16532 5322 16544
rect 5629 16541 5641 16544
rect 5675 16572 5687 16575
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 5675 16544 5825 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 5997 16575 6055 16581
rect 5997 16541 6009 16575
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 5353 16507 5411 16513
rect 5353 16504 5365 16507
rect 4396 16476 5365 16504
rect 4396 16464 4402 16476
rect 5353 16473 5365 16476
rect 5399 16473 5411 16507
rect 5353 16467 5411 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 4246 16436 4252 16448
rect 3283 16408 4252 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 4982 16396 4988 16448
rect 5040 16396 5046 16448
rect 5626 16396 5632 16448
rect 5684 16436 5690 16448
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5684 16408 5917 16436
rect 5684 16396 5690 16408
rect 5905 16405 5917 16408
rect 5951 16405 5963 16439
rect 6012 16436 6040 16535
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 9272 16544 12173 16572
rect 9272 16532 9278 16544
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 6086 16464 6092 16516
rect 6144 16504 6150 16516
rect 7101 16507 7159 16513
rect 7101 16504 7113 16507
rect 6144 16476 7113 16504
rect 6144 16464 6150 16476
rect 7101 16473 7113 16476
rect 7147 16473 7159 16507
rect 7101 16467 7159 16473
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 8294 16504 8300 16516
rect 7800 16476 8300 16504
rect 7800 16464 7806 16476
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 12069 16507 12127 16513
rect 12069 16473 12081 16507
rect 12115 16473 12127 16507
rect 12069 16467 12127 16473
rect 6270 16436 6276 16448
rect 6012 16408 6276 16436
rect 5905 16399 5963 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11848 16408 11897 16436
rect 11848 16396 11854 16408
rect 11885 16405 11897 16408
rect 11931 16436 11943 16439
rect 12084 16436 12112 16467
rect 11931 16408 12112 16436
rect 12268 16436 12296 16612
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 13170 16640 13176 16652
rect 12391 16612 13176 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 14182 16600 14188 16652
rect 14240 16600 14246 16652
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12897 16575 12955 16581
rect 12897 16572 12909 16575
rect 12492 16544 12909 16572
rect 12492 16532 12498 16544
rect 12897 16541 12909 16544
rect 12943 16541 12955 16575
rect 12897 16535 12955 16541
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 15654 16572 15660 16584
rect 14415 16544 15660 16572
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 12526 16464 12532 16516
rect 12584 16464 12590 16516
rect 13280 16504 13308 16535
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 13725 16507 13783 16513
rect 13725 16504 13737 16507
rect 13280 16476 13737 16504
rect 13280 16436 13308 16476
rect 13725 16473 13737 16476
rect 13771 16473 13783 16507
rect 13725 16467 13783 16473
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 12268 16408 13308 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 14568 16436 14596 16467
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15197 16507 15255 16513
rect 15197 16504 15209 16507
rect 14884 16476 15209 16504
rect 14884 16464 14890 16476
rect 15197 16473 15209 16476
rect 15243 16473 15255 16507
rect 15197 16467 15255 16473
rect 14918 16436 14924 16448
rect 14568 16408 14924 16436
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 1104 16346 18860 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 18860 16346
rect 1104 16272 18860 16294
rect 8202 16232 8208 16244
rect 4172 16204 8208 16232
rect 4172 16173 4200 16204
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 10744 16204 14841 16232
rect 10744 16192 10750 16204
rect 14829 16201 14841 16204
rect 14875 16232 14887 16235
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 14875 16204 15117 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 15105 16195 15163 16201
rect 4157 16167 4215 16173
rect 4157 16133 4169 16167
rect 4203 16133 4215 16167
rect 5810 16164 5816 16176
rect 5474 16136 5816 16164
rect 4157 16127 4215 16133
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 5902 16124 5908 16176
rect 5960 16124 5966 16176
rect 5994 16124 6000 16176
rect 6052 16164 6058 16176
rect 8110 16164 8116 16176
rect 6052 16136 8116 16164
rect 6052 16124 6058 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 15194 16164 15200 16176
rect 12558 16136 15200 16164
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 14884 16068 15025 16096
rect 14884 16056 14890 16068
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15289 16099 15347 16105
rect 15289 16065 15301 16099
rect 15335 16096 15347 16099
rect 15470 16096 15476 16108
rect 15335 16068 15476 16096
rect 15335 16065 15347 16068
rect 15289 16059 15347 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 6178 15988 6184 16040
rect 6236 15988 6242 16040
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 11238 16028 11244 16040
rect 6420 16000 11244 16028
rect 6420 15988 6426 16000
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 12986 15988 12992 16040
rect 13044 15988 13050 16040
rect 17402 16028 17408 16040
rect 13188 16000 17408 16028
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3786 15892 3792 15904
rect 3099 15864 3792 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 5868 15864 11529 15892
rect 5868 15852 5874 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 13188 15892 13216 16000
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 14752 15932 15485 15960
rect 14752 15904 14780 15932
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 15473 15923 15531 15929
rect 12676 15864 13216 15892
rect 14001 15895 14059 15901
rect 12676 15852 12682 15864
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14458 15892 14464 15904
rect 14047 15864 14464 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 14553 15895 14611 15901
rect 14553 15861 14565 15895
rect 14599 15892 14611 15895
rect 14734 15892 14740 15904
rect 14599 15864 14740 15892
rect 14599 15861 14611 15864
rect 14553 15855 14611 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 15378 15852 15384 15904
rect 15436 15852 15442 15904
rect 15749 15895 15807 15901
rect 15749 15861 15761 15895
rect 15795 15892 15807 15895
rect 16298 15892 16304 15904
rect 15795 15864 16304 15892
rect 15795 15861 15807 15864
rect 15749 15855 15807 15861
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 1104 15802 18860 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 18860 15802
rect 1104 15728 18860 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 6362 15688 6368 15700
rect 3651 15660 6368 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 3878 15580 3884 15632
rect 3936 15620 3942 15632
rect 7653 15623 7711 15629
rect 7653 15620 7665 15623
rect 3936 15592 7665 15620
rect 3936 15580 3942 15592
rect 7653 15589 7665 15592
rect 7699 15589 7711 15623
rect 7852 15620 7880 15651
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8754 15688 8760 15700
rect 8260 15660 8760 15688
rect 8260 15648 8266 15660
rect 8754 15648 8760 15660
rect 8812 15688 8818 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 8812 15660 10057 15688
rect 8812 15648 8818 15660
rect 10045 15657 10057 15660
rect 10091 15688 10103 15691
rect 10091 15660 10765 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 7852 15592 9520 15620
rect 7653 15583 7711 15589
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 2498 15552 2504 15564
rect 1903 15524 2504 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 2498 15512 2504 15524
rect 2556 15552 2562 15564
rect 6178 15552 6184 15564
rect 2556 15524 6184 15552
rect 2556 15512 2562 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 6362 15552 6368 15564
rect 6319 15524 6368 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 6362 15512 6368 15524
rect 6420 15552 6426 15564
rect 6638 15552 6644 15564
rect 6420 15524 6644 15552
rect 6420 15512 6426 15524
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7340 15524 7481 15552
rect 7340 15512 7346 15524
rect 7469 15521 7481 15524
rect 7515 15552 7527 15555
rect 8018 15552 8024 15564
rect 7515 15524 8024 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 1578 15484 1584 15496
rect 1443 15456 1584 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 4430 15484 4436 15496
rect 3266 15456 4436 15484
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4672 15456 5273 15484
rect 4672 15444 4678 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5442 15444 5448 15496
rect 5500 15444 5506 15496
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 9492 15484 9520 15592
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 10410 15620 10416 15632
rect 9640 15592 10416 15620
rect 9640 15580 9646 15592
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 10737 15552 10765 15660
rect 11238 15648 11244 15700
rect 11296 15648 11302 15700
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13228 15660 14105 15688
rect 13228 15648 13234 15660
rect 14093 15657 14105 15660
rect 14139 15688 14151 15691
rect 15838 15688 15844 15700
rect 14139 15660 15844 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 11517 15623 11575 15629
rect 11517 15589 11529 15623
rect 11563 15620 11575 15623
rect 12618 15620 12624 15632
rect 11563 15592 12624 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 16574 15620 16580 15632
rect 13412 15592 16580 15620
rect 13412 15580 13418 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 10737 15524 10824 15552
rect 10318 15484 10324 15496
rect 5859 15456 9444 15484
rect 9492 15456 10324 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 2130 15376 2136 15428
rect 2188 15416 2194 15428
rect 3973 15419 4031 15425
rect 3973 15416 3985 15419
rect 2188 15388 2544 15416
rect 2188 15376 2194 15388
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 2406 15348 2412 15360
rect 1627 15320 2412 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2516 15348 2544 15388
rect 3436 15388 3985 15416
rect 3436 15348 3464 15388
rect 3973 15385 3985 15388
rect 4019 15385 4031 15419
rect 3973 15379 4031 15385
rect 4525 15419 4583 15425
rect 4525 15385 4537 15419
rect 4571 15385 4583 15419
rect 4525 15379 4583 15385
rect 2516 15320 3464 15348
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 4341 15351 4399 15357
rect 4341 15348 4353 15351
rect 4120 15320 4353 15348
rect 4120 15308 4126 15320
rect 4341 15317 4353 15320
rect 4387 15348 4399 15351
rect 4540 15348 4568 15379
rect 4706 15376 4712 15428
rect 4764 15376 4770 15428
rect 4890 15376 4896 15428
rect 4948 15376 4954 15428
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15416 5687 15419
rect 5994 15416 6000 15428
rect 5675 15388 6000 15416
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 7834 15425 7840 15428
rect 7193 15419 7251 15425
rect 7193 15385 7205 15419
rect 7239 15416 7251 15419
rect 7821 15419 7840 15425
rect 7821 15416 7833 15419
rect 7239 15388 7833 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 7821 15385 7833 15388
rect 7821 15379 7840 15385
rect 7834 15376 7840 15379
rect 7892 15376 7898 15428
rect 8018 15376 8024 15428
rect 8076 15376 8082 15428
rect 9416 15416 9444 15456
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10796 15493 10824 15524
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 11112 15524 12173 15552
rect 11112 15512 11118 15524
rect 11716 15496 11744 15524
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 15286 15552 15292 15564
rect 12161 15515 12219 15521
rect 13096 15524 15292 15552
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 10781 15487 10839 15493
rect 10643 15456 10677 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10781 15453 10793 15487
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 9582 15416 9588 15428
rect 9416 15388 9588 15416
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 10505 15419 10563 15425
rect 10505 15385 10517 15419
rect 10551 15416 10563 15419
rect 10612 15416 10640 15447
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11296 15456 11437 15484
rect 11296 15444 11302 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15484 11851 15487
rect 13096 15484 13124 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 11839 15456 13124 15484
rect 14369 15487 14427 15493
rect 11839 15453 11851 15456
rect 11793 15447 11851 15453
rect 14369 15453 14381 15487
rect 14415 15484 14427 15487
rect 14458 15484 14464 15496
rect 14415 15456 14464 15484
rect 14415 15453 14427 15456
rect 14369 15447 14427 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 13630 15416 13636 15428
rect 10551 15388 13636 15416
rect 10551 15385 10563 15388
rect 10505 15379 10563 15385
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 13817 15419 13875 15425
rect 13817 15385 13829 15419
rect 13863 15416 13875 15419
rect 14645 15419 14703 15425
rect 13863 15388 14320 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 14292 15360 14320 15388
rect 14645 15385 14657 15419
rect 14691 15416 14703 15419
rect 15654 15416 15660 15428
rect 14691 15388 15660 15416
rect 14691 15385 14703 15388
rect 14645 15379 14703 15385
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 4387 15320 4568 15348
rect 5077 15351 5135 15357
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 5258 15348 5264 15360
rect 5123 15320 5264 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15348 5411 15351
rect 6641 15351 6699 15357
rect 6641 15348 6653 15351
rect 5399 15320 6653 15348
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 6641 15317 6653 15320
rect 6687 15348 6699 15351
rect 8478 15348 8484 15360
rect 6687 15320 8484 15348
rect 6687 15317 6699 15320
rect 6641 15311 6699 15317
rect 8478 15308 8484 15320
rect 8536 15348 8542 15360
rect 9398 15348 9404 15360
rect 8536 15320 9404 15348
rect 8536 15308 8542 15320
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 10594 15308 10600 15360
rect 10652 15308 10658 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14461 15351 14519 15357
rect 14461 15317 14473 15351
rect 14507 15348 14519 15351
rect 15010 15348 15016 15360
rect 14507 15320 15016 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15562 15348 15568 15360
rect 15335 15320 15568 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 18506 15308 18512 15360
rect 18564 15308 18570 15360
rect 1104 15258 18860 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 18860 15258
rect 1104 15184 18860 15206
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 13722 15144 13728 15156
rect 10827 15116 13728 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13998 15153 14004 15156
rect 13985 15147 14004 15153
rect 13985 15113 13997 15147
rect 13985 15107 14004 15113
rect 13998 15104 14004 15107
rect 14056 15104 14062 15156
rect 15194 15104 15200 15156
rect 15252 15104 15258 15156
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 15304 15116 15761 15144
rect 1578 15036 1584 15088
rect 1636 15036 1642 15088
rect 5169 15079 5227 15085
rect 5169 15045 5181 15079
rect 5215 15076 5227 15079
rect 5813 15079 5871 15085
rect 5813 15076 5825 15079
rect 5215 15048 5825 15076
rect 5215 15045 5227 15048
rect 5169 15039 5227 15045
rect 5813 15045 5825 15048
rect 5859 15076 5871 15079
rect 6086 15076 6092 15088
rect 5859 15048 6092 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6086 15036 6092 15048
rect 6144 15036 6150 15088
rect 6454 15036 6460 15088
rect 6512 15076 6518 15088
rect 9306 15076 9312 15088
rect 6512 15048 9312 15076
rect 6512 15036 6518 15048
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 9490 15085 9496 15088
rect 9477 15079 9496 15085
rect 9477 15045 9489 15079
rect 9477 15039 9496 15045
rect 9490 15036 9496 15039
rect 9548 15036 9554 15088
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 10134 15076 10140 15088
rect 9723 15048 10140 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 14182 15036 14188 15088
rect 14240 15036 14246 15088
rect 14826 15036 14832 15088
rect 14884 15076 14890 15088
rect 15304 15076 15332 15116
rect 15749 15113 15761 15116
rect 15795 15113 15807 15147
rect 15749 15107 15807 15113
rect 14884 15048 15332 15076
rect 14884 15036 14890 15048
rect 15562 15036 15568 15088
rect 15620 15076 15626 15088
rect 15620 15048 15884 15076
rect 15620 15036 15626 15048
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 5718 15008 5724 15020
rect 5675 14980 5724 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 14977 5963 15011
rect 6104 15008 6132 15036
rect 15856 15017 15884 15048
rect 10045 15011 10103 15017
rect 10045 15008 10057 15011
rect 6104 14980 10057 15008
rect 5905 14971 5963 14977
rect 10045 14977 10057 14980
rect 10091 15008 10103 15011
rect 10722 15011 10780 15017
rect 10722 15008 10734 15011
rect 10091 14980 10734 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10722 14977 10734 14980
rect 10768 14977 10780 15011
rect 10722 14971 10780 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 15059 14980 15301 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15289 14977 15301 14980
rect 15335 15008 15347 15011
rect 15841 15011 15899 15017
rect 15335 14980 15516 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 5920 14940 5948 14971
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 4080 14912 6653 14940
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 2372 14776 2421 14804
rect 2372 14764 2378 14776
rect 2409 14773 2421 14776
rect 2455 14804 2467 14807
rect 4080 14804 4108 14912
rect 6641 14909 6653 14912
rect 6687 14940 6699 14943
rect 10318 14940 10324 14952
rect 6687 14912 10324 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10594 14940 10600 14952
rect 10551 14912 10600 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 10928 14912 11253 14940
rect 10928 14900 10934 14912
rect 11241 14909 11253 14912
rect 11287 14940 11299 14943
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11287 14912 11713 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 15381 14943 15439 14949
rect 11701 14903 11759 14909
rect 13556 14912 14688 14940
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 5629 14875 5687 14881
rect 5629 14872 5641 14875
rect 4212 14844 5641 14872
rect 4212 14832 4218 14844
rect 5629 14841 5641 14844
rect 5675 14841 5687 14875
rect 5629 14835 5687 14841
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6362 14872 6368 14884
rect 5776 14844 6368 14872
rect 5776 14832 5782 14844
rect 6362 14832 6368 14844
rect 6420 14872 6426 14884
rect 13556 14872 13584 14912
rect 6420 14844 13584 14872
rect 13648 14844 14044 14872
rect 6420 14832 6426 14844
rect 2455 14776 4108 14804
rect 5537 14807 5595 14813
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 5736 14804 5764 14832
rect 5583 14776 5764 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 8386 14804 8392 14816
rect 6236 14776 8392 14804
rect 6236 14764 6242 14776
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 9180 14776 9321 14804
rect 9180 14764 9186 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9309 14767 9367 14773
rect 9490 14764 9496 14816
rect 9548 14764 9554 14816
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 10686 14764 10692 14816
rect 10744 14804 10750 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 10744 14776 11161 14804
rect 10744 14764 10750 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 13648 14813 13676 14844
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 12400 14776 13645 14804
rect 12400 14764 12406 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14804 13875 14807
rect 13906 14804 13912 14816
rect 13863 14776 13912 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14016 14813 14044 14844
rect 14660 14813 14688 14912
rect 15381 14909 15393 14943
rect 15427 14909 15439 14943
rect 15488 14940 15516 14980
rect 15841 14977 15853 15011
rect 15887 14977 15899 15011
rect 15841 14971 15899 14977
rect 16482 14940 16488 14952
rect 15488 14912 16488 14940
rect 15381 14903 15439 14909
rect 15396 14872 15424 14903
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16022 14872 16028 14884
rect 15396 14844 16028 14872
rect 16022 14832 16028 14844
rect 16080 14832 16086 14884
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14773 14059 14807
rect 14001 14767 14059 14773
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 14826 14804 14832 14816
rect 14691 14776 14832 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 18598 14804 18604 14816
rect 15611 14776 18604 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 1104 14714 18860 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 18860 14714
rect 1104 14640 18860 14662
rect 2225 14603 2283 14609
rect 2225 14569 2237 14603
rect 2271 14569 2283 14603
rect 2225 14563 2283 14569
rect 2240 14532 2268 14563
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3568 14572 4169 14600
rect 3568 14560 3574 14572
rect 4157 14569 4169 14572
rect 4203 14600 4215 14603
rect 4338 14600 4344 14612
rect 4203 14572 4344 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 6454 14600 6460 14612
rect 4724 14572 6460 14600
rect 2593 14535 2651 14541
rect 2593 14532 2605 14535
rect 2240 14504 2605 14532
rect 2593 14501 2605 14504
rect 2639 14532 2651 14535
rect 4724 14532 4752 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 7374 14600 7380 14612
rect 6696 14572 7380 14600
rect 6696 14560 6702 14572
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 7800 14572 8340 14600
rect 7800 14560 7806 14572
rect 2639 14504 4752 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 5718 14492 5724 14544
rect 5776 14532 5782 14544
rect 5994 14532 6000 14544
rect 5776 14504 6000 14532
rect 5776 14492 5782 14504
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 8312 14532 8340 14572
rect 9398 14560 9404 14612
rect 9456 14600 9462 14612
rect 9769 14603 9827 14609
rect 9769 14600 9781 14603
rect 9456 14572 9781 14600
rect 9456 14560 9462 14572
rect 9769 14569 9781 14572
rect 9815 14569 9827 14603
rect 13354 14600 13360 14612
rect 9769 14563 9827 14569
rect 9876 14572 13360 14600
rect 9876 14532 9904 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 8312 14504 9904 14532
rect 12621 14535 12679 14541
rect 12621 14501 12633 14535
rect 12667 14532 12679 14535
rect 12667 14504 16160 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 2148 14436 3433 14464
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 2148 14405 2176 14436
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 5074 14424 5080 14476
rect 5132 14424 5138 14476
rect 5166 14424 5172 14476
rect 5224 14464 5230 14476
rect 7466 14464 7472 14476
rect 5224 14436 7472 14464
rect 5224 14424 5230 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 11974 14464 11980 14476
rect 8168 14436 11980 14464
rect 8168 14424 8174 14436
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12124 14436 12357 14464
rect 12124 14424 12130 14436
rect 12345 14433 12357 14436
rect 12391 14464 12403 14467
rect 12391 14436 12756 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 1728 14368 2145 14396
rect 1728 14356 1734 14368
rect 2133 14365 2145 14368
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2314 14396 2320 14408
rect 2271 14368 2320 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2685 14399 2743 14405
rect 2685 14396 2697 14399
rect 2464 14368 2697 14396
rect 2464 14356 2470 14368
rect 2685 14365 2697 14368
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3786 14396 3792 14408
rect 3007 14368 3792 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5092 14396 5120 14424
rect 4948 14368 6132 14396
rect 4948 14356 4954 14368
rect 4525 14331 4583 14337
rect 4525 14297 4537 14331
rect 4571 14328 4583 14331
rect 5074 14328 5080 14340
rect 4571 14300 5080 14328
rect 4571 14297 4583 14300
rect 4525 14291 4583 14297
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 1857 14263 1915 14269
rect 1857 14229 1869 14263
rect 1903 14260 1915 14263
rect 2314 14260 2320 14272
rect 1903 14232 2320 14260
rect 1903 14229 1915 14232
rect 1857 14223 1915 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 5994 14220 6000 14272
rect 6052 14220 6058 14272
rect 6104 14260 6132 14368
rect 8386 14356 8392 14408
rect 8444 14356 8450 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12728 14405 12756 14436
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 14366 14464 14372 14476
rect 13596 14436 14372 14464
rect 13596 14424 13602 14436
rect 14366 14424 14372 14436
rect 14424 14464 14430 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14424 14436 15485 14464
rect 14424 14424 14430 14436
rect 15473 14433 15485 14436
rect 15519 14464 15531 14467
rect 15746 14464 15752 14476
rect 15519 14436 15752 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 16132 14464 16160 14504
rect 17310 14492 17316 14544
rect 17368 14532 17374 14544
rect 18325 14535 18383 14541
rect 18325 14532 18337 14535
rect 17368 14504 18337 14532
rect 17368 14492 17374 14504
rect 18325 14501 18337 14504
rect 18371 14501 18383 14535
rect 18325 14495 18383 14501
rect 17494 14464 17500 14476
rect 16132 14436 17500 14464
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 12492 14368 12541 14396
rect 12492 14356 12498 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15160 14368 16037 14396
rect 15160 14356 15166 14368
rect 16025 14365 16037 14368
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18874 14396 18880 14408
rect 18555 14368 18880 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 7682 14300 8064 14328
rect 7742 14260 7748 14272
rect 6104 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8036 14260 8064 14300
rect 8110 14288 8116 14340
rect 8168 14288 8174 14340
rect 11238 14328 11244 14340
rect 8220 14300 11244 14328
rect 8220 14260 8248 14300
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 16301 14331 16359 14337
rect 16301 14328 16313 14331
rect 15344 14300 16313 14328
rect 15344 14288 15350 14300
rect 16301 14297 16313 14300
rect 16347 14297 16359 14331
rect 16301 14291 16359 14297
rect 16850 14288 16856 14340
rect 16908 14288 16914 14340
rect 8036 14232 8248 14260
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 16206 14260 16212 14272
rect 11388 14232 16212 14260
rect 11388 14220 11394 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 17773 14263 17831 14269
rect 17773 14260 17785 14263
rect 16448 14232 17785 14260
rect 16448 14220 16454 14232
rect 17773 14229 17785 14232
rect 17819 14229 17831 14263
rect 17773 14223 17831 14229
rect 18230 14220 18236 14272
rect 18288 14220 18294 14272
rect 1104 14170 18860 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 18860 14170
rect 1104 14096 18860 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4890 14056 4896 14068
rect 4203 14028 4896 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 3881 13991 3939 13997
rect 3881 13957 3893 13991
rect 3927 13988 3939 13991
rect 4062 13988 4068 14000
rect 3927 13960 4068 13988
rect 3927 13957 3939 13960
rect 3881 13951 3939 13957
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 4172 13920 4200 14019
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 6565 14059 6623 14065
rect 6565 14056 6577 14059
rect 5040 14028 6577 14056
rect 5040 14016 5046 14028
rect 6565 14025 6577 14028
rect 6611 14025 6623 14059
rect 6565 14019 6623 14025
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 7282 14056 7288 14068
rect 6840 14028 7288 14056
rect 5166 13948 5172 14000
rect 5224 13948 5230 14000
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 5629 13991 5687 13997
rect 5629 13988 5641 13991
rect 5592 13960 5641 13988
rect 5592 13948 5598 13960
rect 5629 13957 5641 13960
rect 5675 13988 5687 13991
rect 5994 13988 6000 14000
rect 5675 13960 6000 13988
rect 5675 13957 5687 13960
rect 5629 13951 5687 13957
rect 5994 13948 6000 13960
rect 6052 13948 6058 14000
rect 6365 13991 6423 13997
rect 6365 13957 6377 13991
rect 6411 13988 6423 13991
rect 6454 13988 6460 14000
rect 6411 13960 6460 13988
rect 6411 13957 6423 13960
rect 6365 13951 6423 13957
rect 6454 13948 6460 13960
rect 6512 13988 6518 14000
rect 6840 13988 6868 14028
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7340 14028 8401 14056
rect 7340 14016 7346 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 8720 14028 11529 14056
rect 8720 14016 8726 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 12032 14028 13369 14056
rect 12032 14016 12038 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 16264 14028 17417 14056
rect 16264 14016 16270 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 8113 13991 8171 13997
rect 8113 13988 8125 13991
rect 6512 13960 6868 13988
rect 7024 13960 8125 13988
rect 6512 13948 6518 13960
rect 4019 13892 4200 13920
rect 5905 13923 5963 13929
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 6178 13920 6184 13932
rect 5951 13892 6184 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 2406 13812 2412 13864
rect 2464 13852 2470 13864
rect 2590 13852 2596 13864
rect 2464 13824 2596 13852
rect 2464 13812 2470 13824
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3804 13852 3832 13883
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 7024 13929 7052 13960
rect 8113 13957 8125 13960
rect 8159 13988 8171 13991
rect 9398 13988 9404 14000
rect 8159 13960 9404 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 11669 13991 11727 13997
rect 11669 13988 11681 13991
rect 11480 13960 11681 13988
rect 11480 13948 11486 13960
rect 11669 13957 11681 13960
rect 11715 13957 11727 13991
rect 11669 13951 11727 13957
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 12342 13988 12348 14000
rect 11931 13960 12348 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 13320 13960 13860 13988
rect 13320 13948 13326 13960
rect 13832 13932 13860 13960
rect 14090 13948 14096 14000
rect 14148 13948 14154 14000
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 15804 13960 15884 13988
rect 15804 13948 15810 13960
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13920 7251 13923
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7239 13892 7757 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7745 13889 7757 13892
rect 7791 13920 7803 13923
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 7791 13892 10241 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 10229 13889 10241 13892
rect 10275 13920 10287 13923
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10275 13892 10517 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10505 13889 10517 13892
rect 10551 13920 10563 13923
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 10551 13910 12296 13920
rect 12452 13910 13093 13920
rect 10551 13892 13093 13910
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 12268 13882 12480 13892
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 13127 13892 13461 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13449 13889 13461 13892
rect 13495 13920 13507 13923
rect 13538 13920 13544 13932
rect 13495 13892 13544 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 15856 13929 15884 13960
rect 15841 13923 15899 13929
rect 15841 13889 15853 13923
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16114 13880 16120 13932
rect 16172 13880 16178 13932
rect 17420 13920 17448 14019
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 18012 14028 18061 14056
rect 18012 14016 18018 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 17932 13923 17990 13929
rect 17932 13920 17944 13923
rect 17420 13892 17944 13920
rect 17932 13889 17944 13892
rect 17978 13889 17990 13923
rect 17932 13883 17990 13889
rect 5074 13852 5080 13864
rect 3804 13824 5080 13852
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 5224 13824 6929 13852
rect 5224 13812 5230 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 7466 13852 7472 13864
rect 7331 13824 7472 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 8996 13824 10149 13852
rect 8996 13812 9002 13824
rect 10137 13821 10149 13824
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 15565 13855 15623 13861
rect 10468 13824 15148 13852
rect 10468 13812 10474 13824
rect 12710 13784 12716 13796
rect 5828 13756 10180 13784
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5828 13716 5856 13756
rect 10152 13728 10180 13756
rect 11716 13756 12716 13784
rect 4948 13688 5856 13716
rect 4948 13676 4954 13688
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6454 13716 6460 13728
rect 6052 13688 6460 13716
rect 6052 13676 6058 13688
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 6546 13676 6552 13728
rect 6604 13676 6610 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 9674 13716 9680 13728
rect 6696 13688 9680 13716
rect 6696 13676 6702 13688
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 11716 13725 11744 13756
rect 12710 13744 12716 13756
rect 12768 13744 12774 13796
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13262 13784 13268 13796
rect 12860 13756 13268 13784
rect 12860 13744 12866 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 15120 13784 15148 13824
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 15654 13852 15660 13864
rect 15611 13824 15660 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17310 13852 17316 13864
rect 17175 13824 17316 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17310 13812 17316 13824
rect 17368 13852 17374 13864
rect 17368 13824 17816 13852
rect 17368 13812 17374 13824
rect 17788 13784 17816 13824
rect 18138 13812 18144 13864
rect 18196 13812 18202 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18248 13824 18429 13852
rect 18248 13784 18276 13824
rect 18417 13821 18429 13824
rect 18463 13821 18475 13855
rect 18417 13815 18475 13821
rect 15120 13756 16436 13784
rect 17788 13756 18276 13784
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13685 11759 13719
rect 11701 13679 11759 13685
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12342 13716 12348 13728
rect 12299 13688 12348 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 16298 13716 16304 13728
rect 12952 13688 16304 13716
rect 12952 13676 12958 13688
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 16408 13716 16436 13756
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 16408 13688 17785 13716
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 1104 13626 18860 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 18860 13626
rect 1104 13552 18860 13574
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 4982 13512 4988 13524
rect 4488 13484 4988 13512
rect 4488 13472 4494 13484
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 5500 13484 8125 13512
rect 5500 13472 5506 13484
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 4890 13376 4896 13388
rect 4755 13348 4896 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 6178 13336 6184 13388
rect 6236 13376 6242 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6236 13348 6469 13376
rect 6236 13336 6242 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 3878 13268 3884 13320
rect 3936 13268 3942 13320
rect 4430 13268 4436 13320
rect 4488 13268 4494 13320
rect 6748 13317 6776 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 12894 13512 12900 13524
rect 8113 13475 8171 13481
rect 8220 13484 12900 13512
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 8220 13444 8248 13484
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 16114 13512 16120 13524
rect 13004 13484 16120 13512
rect 6880 13416 8248 13444
rect 6880 13404 6886 13416
rect 8110 13376 8116 13388
rect 6932 13348 8116 13376
rect 6932 13317 6960 13348
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10376 13348 11284 13376
rect 10376 13336 10382 13348
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13277 6791 13311
rect 6733 13271 6791 13277
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13277 7343 13311
rect 7285 13271 7343 13277
rect 5166 13200 5172 13252
rect 5224 13200 5230 13252
rect 6181 13243 6239 13249
rect 6181 13209 6193 13243
rect 6227 13240 6239 13243
rect 6454 13240 6460 13252
rect 6227 13212 6460 13240
rect 6227 13209 6239 13212
rect 6181 13203 6239 13209
rect 6454 13200 6460 13212
rect 6512 13200 6518 13252
rect 7300 13240 7328 13271
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7432 13280 7481 13308
rect 7432 13268 7438 13280
rect 7469 13277 7481 13280
rect 7515 13308 7527 13311
rect 8481 13311 8539 13317
rect 8481 13308 8493 13311
rect 7515 13280 8493 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 8481 13277 8493 13280
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 10008 13280 10241 13308
rect 10008 13268 10014 13280
rect 10229 13277 10241 13280
rect 10275 13308 10287 13311
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10275 13280 10609 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 7837 13243 7895 13249
rect 7837 13240 7849 13243
rect 7300 13212 7849 13240
rect 7837 13209 7849 13212
rect 7883 13240 7895 13243
rect 8202 13240 8208 13252
rect 7883 13212 8208 13240
rect 7883 13209 7895 13212
rect 7837 13203 7895 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 10505 13243 10563 13249
rect 10505 13240 10517 13243
rect 9088 13212 10517 13240
rect 9088 13200 9094 13212
rect 10505 13209 10517 13212
rect 10551 13209 10563 13243
rect 11256 13240 11284 13348
rect 13004 13317 13032 13484
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17460 13484 17540 13512
rect 17460 13472 17466 13484
rect 17512 13444 17540 13484
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 17644 13484 17693 13512
rect 17644 13472 17650 13484
rect 17681 13481 17693 13484
rect 17727 13512 17739 13515
rect 17862 13512 17868 13524
rect 17727 13484 17868 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 18012 13484 18061 13512
rect 18012 13472 18018 13484
rect 18049 13481 18061 13484
rect 18095 13512 18107 13515
rect 18138 13512 18144 13524
rect 18095 13484 18144 13512
rect 18095 13481 18107 13484
rect 18049 13475 18107 13481
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 17512 13416 18184 13444
rect 18156 13388 18184 13416
rect 13722 13376 13728 13388
rect 13096 13348 13728 13376
rect 13096 13317 13124 13348
rect 13722 13336 13728 13348
rect 13780 13376 13786 13388
rect 14642 13376 14648 13388
rect 13780 13348 14648 13376
rect 13780 13336 13786 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 18138 13336 18144 13388
rect 18196 13336 18202 13388
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13188 13240 13216 13271
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 15120 13308 15148 13336
rect 15286 13308 15292 13320
rect 13872 13280 15292 13308
rect 13872 13268 13878 13280
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 13449 13243 13507 13249
rect 13449 13240 13461 13243
rect 11256 13212 13461 13240
rect 10505 13203 10563 13209
rect 13449 13209 13461 13212
rect 13495 13209 13507 13243
rect 13449 13203 13507 13209
rect 3602 13132 3608 13184
rect 3660 13172 3666 13184
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 3660 13144 4077 13172
rect 3660 13132 3666 13144
rect 4065 13141 4077 13144
rect 4111 13141 4123 13175
rect 4065 13135 4123 13141
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 6638 13172 6644 13184
rect 4663 13144 6644 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 6788 13144 6837 13172
rect 6788 13132 6794 13144
rect 6825 13141 6837 13144
rect 6871 13141 6883 13175
rect 6825 13135 6883 13141
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 6972 13144 7389 13172
rect 6972 13132 6978 13144
rect 7377 13141 7389 13144
rect 7423 13141 7435 13175
rect 7377 13135 7435 13141
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 12802 13172 12808 13184
rect 7616 13144 12808 13172
rect 7616 13132 7622 13144
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13464 13172 13492 13203
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 13688 13212 15577 13240
rect 13688 13200 13694 13212
rect 15565 13209 15577 13212
rect 15611 13209 15623 13243
rect 15565 13203 15623 13209
rect 16574 13200 16580 13252
rect 16632 13200 16638 13252
rect 17313 13243 17371 13249
rect 17313 13209 17325 13243
rect 17359 13209 17371 13243
rect 17313 13203 17371 13209
rect 17328 13172 17356 13203
rect 13464 13144 17356 13172
rect 18506 13132 18512 13184
rect 18564 13132 18570 13184
rect 1104 13082 18860 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 18860 13082
rect 1104 13008 18860 13030
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 6822 12968 6828 12980
rect 2823 12940 6828 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2884 12841 2912 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 10042 12968 10048 12980
rect 7836 12940 10048 12968
rect 3694 12860 3700 12912
rect 3752 12860 3758 12912
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 6236 12872 6469 12900
rect 6236 12860 6242 12872
rect 6457 12869 6469 12872
rect 6503 12900 6515 12903
rect 7742 12900 7748 12912
rect 6503 12872 7748 12900
rect 6503 12869 6515 12872
rect 6457 12863 6515 12869
rect 7742 12860 7748 12872
rect 7800 12860 7806 12912
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3510 12832 3516 12844
rect 3016 12804 3516 12832
rect 3016 12792 3022 12804
rect 3510 12792 3516 12804
rect 3568 12832 3574 12844
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3568 12804 3617 12832
rect 3568 12792 3574 12804
rect 3605 12801 3617 12804
rect 3651 12832 3663 12835
rect 3786 12832 3792 12844
rect 3651 12804 3792 12832
rect 3651 12801 3663 12804
rect 3605 12795 3663 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6932 12804 7021 12832
rect 1762 12724 1768 12776
rect 1820 12764 1826 12776
rect 6932 12764 6960 12804
rect 7009 12801 7021 12804
rect 7055 12832 7067 12835
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7055 12804 7573 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7561 12801 7573 12804
rect 7607 12832 7619 12835
rect 7836 12832 7864 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10428 12940 11468 12968
rect 8570 12860 8576 12912
rect 8628 12860 8634 12912
rect 10428 12841 10456 12940
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 11117 12903 11175 12909
rect 11117 12900 11129 12903
rect 11020 12872 11129 12900
rect 11020 12860 11026 12872
rect 11117 12869 11129 12872
rect 11163 12869 11175 12903
rect 11117 12863 11175 12869
rect 11333 12903 11391 12909
rect 11333 12869 11345 12903
rect 11379 12869 11391 12903
rect 11440 12900 11468 12940
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 11572 12940 18429 12968
rect 11572 12928 11578 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 15562 12900 15568 12912
rect 11440 12872 15568 12900
rect 11333 12863 11391 12869
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 7607 12804 7864 12832
rect 10244 12804 10425 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 1820 12736 6960 12764
rect 7837 12767 7895 12773
rect 1820 12724 1826 12736
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7837 12727 7895 12733
rect 7944 12736 8125 12764
rect 3050 12656 3056 12708
rect 3108 12656 3114 12708
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 5994 12696 6000 12708
rect 4120 12668 6000 12696
rect 4120 12656 4126 12668
rect 5994 12656 6000 12668
rect 6052 12696 6058 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 6052 12668 7205 12696
rect 6052 12656 6058 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 7852 12696 7880 12727
rect 7800 12668 7880 12696
rect 7800 12656 7806 12668
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 6362 12628 6368 12640
rect 5592 12600 6368 12628
rect 5592 12588 5598 12600
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 7944 12628 7972 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 10244 12773 10272 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10229 12767 10287 12773
rect 10229 12764 10241 12767
rect 8904 12736 10241 12764
rect 8904 12724 8910 12736
rect 10229 12733 10241 12736
rect 10275 12733 10287 12767
rect 10229 12727 10287 12733
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10520 12764 10548 12795
rect 10376 12736 10548 12764
rect 10704 12764 10732 12795
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11348 12832 11376 12863
rect 15562 12860 15568 12872
rect 15620 12900 15626 12912
rect 15930 12900 15936 12912
rect 15620 12872 15936 12900
rect 15620 12860 15626 12872
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 16574 12900 16580 12912
rect 16356 12872 16580 12900
rect 16356 12860 16362 12872
rect 16574 12860 16580 12872
rect 16632 12860 16638 12912
rect 10836 12804 11376 12832
rect 10836 12792 10842 12804
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11756 12804 12265 12832
rect 11756 12792 11762 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12894 12832 12900 12844
rect 12492 12804 12900 12832
rect 12492 12792 12498 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 15344 12804 16681 12832
rect 15344 12792 15350 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 10704 12736 14596 12764
rect 10376 12724 10382 12736
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 10689 12699 10747 12705
rect 9364 12668 9720 12696
rect 9364 12656 9370 12668
rect 7616 12600 7972 12628
rect 7616 12588 7622 12600
rect 9582 12588 9588 12640
rect 9640 12588 9646 12640
rect 9692 12628 9720 12668
rect 10689 12665 10701 12699
rect 10735 12696 10747 12699
rect 10735 12668 12434 12696
rect 10735 12665 10747 12668
rect 10689 12659 10747 12665
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 9692 12600 10977 12628
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11790 12628 11796 12640
rect 11204 12600 11796 12628
rect 11204 12588 11210 12600
rect 11790 12588 11796 12600
rect 11848 12628 11854 12640
rect 12250 12628 12256 12640
rect 11848 12600 12256 12628
rect 11848 12588 11854 12600
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12406 12628 12434 12668
rect 13906 12656 13912 12708
rect 13964 12656 13970 12708
rect 14568 12696 14596 12736
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 15470 12764 15476 12776
rect 14700 12736 15476 12764
rect 14700 12724 14706 12736
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16264 12736 16957 12764
rect 16264 12724 16270 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 16666 12696 16672 12708
rect 14568 12668 16672 12696
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 17586 12628 17592 12640
rect 12406 12600 17592 12628
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 1104 12538 18860 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 18860 12538
rect 1104 12464 18860 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2222 12424 2228 12436
rect 1995 12396 2228 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2222 12384 2228 12396
rect 2280 12424 2286 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2280 12396 2421 12424
rect 2280 12384 2286 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 3568 12396 5549 12424
rect 3568 12384 3574 12396
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 5537 12387 5595 12393
rect 2593 12359 2651 12365
rect 2593 12325 2605 12359
rect 2639 12356 2651 12359
rect 4430 12356 4436 12368
rect 2639 12328 4436 12356
rect 2639 12325 2651 12328
rect 2593 12319 2651 12325
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 5552 12356 5580 12387
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 7558 12424 7564 12436
rect 6052 12396 7564 12424
rect 6052 12384 6058 12396
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 9214 12424 9220 12436
rect 8076 12396 9220 12424
rect 8076 12384 8082 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 10318 12424 10324 12436
rect 9916 12396 10324 12424
rect 9916 12384 9922 12396
rect 10318 12384 10324 12396
rect 10376 12424 10382 12436
rect 10781 12427 10839 12433
rect 10781 12424 10793 12427
rect 10376 12396 10793 12424
rect 10376 12384 10382 12396
rect 10781 12393 10793 12396
rect 10827 12393 10839 12427
rect 10781 12387 10839 12393
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11882 12424 11888 12436
rect 11756 12396 11888 12424
rect 11756 12384 11762 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 14366 12384 14372 12436
rect 14424 12424 14430 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 14424 12396 14473 12424
rect 14424 12384 14430 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 16850 12424 16856 12436
rect 14783 12396 16856 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17494 12424 17500 12436
rect 17000 12396 17500 12424
rect 17000 12384 17006 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 18230 12424 18236 12436
rect 17644 12396 18236 12424
rect 17644 12384 17650 12396
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 5552 12328 5856 12356
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 3568 12260 5733 12288
rect 3568 12248 3574 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3936 12192 3985 12220
rect 3936 12180 3942 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4338 12220 4344 12232
rect 4111 12192 4344 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5828 12229 5856 12328
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 8294 12356 8300 12368
rect 6696 12328 8300 12356
rect 6696 12316 6702 12328
rect 8294 12316 8300 12328
rect 8352 12356 8358 12368
rect 12158 12356 12164 12368
rect 8352 12328 12164 12356
rect 8352 12316 8358 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 12618 12316 12624 12368
rect 12676 12356 12682 12368
rect 12676 12328 17264 12356
rect 12676 12316 12682 12328
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 6236 12260 6285 12288
rect 6236 12248 6242 12260
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 12250 12288 12256 12300
rect 7524 12260 12256 12288
rect 7524 12248 7530 12260
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 12728 12260 16129 12288
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 10594 12220 10600 12232
rect 5813 12183 5871 12189
rect 6840 12192 10600 12220
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 2271 12124 3004 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2406 12044 2412 12096
rect 2464 12093 2470 12096
rect 2976 12093 3004 12124
rect 3786 12112 3792 12164
rect 3844 12112 3850 12164
rect 6840 12152 6868 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11698 12220 11704 12232
rect 11480 12192 11704 12220
rect 11480 12180 11486 12192
rect 11698 12180 11704 12192
rect 11756 12220 11762 12232
rect 12728 12220 12756 12260
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 11756 12192 12756 12220
rect 11756 12180 11762 12192
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12860 12192 13001 12220
rect 12860 12180 12866 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13262 12220 13268 12232
rect 13219 12192 13268 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13262 12180 13268 12192
rect 13320 12220 13326 12232
rect 13446 12220 13452 12232
rect 13320 12192 13452 12220
rect 13320 12180 13326 12192
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14550 12220 14556 12232
rect 14424 12192 14556 12220
rect 14424 12180 14430 12192
rect 14550 12180 14556 12192
rect 14608 12220 14614 12232
rect 14645 12223 14703 12229
rect 14645 12220 14657 12223
rect 14608 12192 14657 12220
rect 14608 12180 14614 12192
rect 14645 12189 14657 12192
rect 14691 12189 14703 12223
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 14645 12183 14703 12189
rect 15856 12192 16037 12220
rect 4080 12124 6868 12152
rect 2464 12087 2483 12093
rect 2471 12053 2483 12087
rect 2464 12047 2483 12053
rect 2961 12087 3019 12093
rect 2961 12053 2973 12087
rect 3007 12084 3019 12087
rect 3970 12084 3976 12096
rect 3007 12056 3976 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 2464 12044 2470 12047
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4080 12093 4108 12124
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 8021 12155 8079 12161
rect 8021 12152 8033 12155
rect 6972 12124 8033 12152
rect 6972 12112 6978 12124
rect 8021 12121 8033 12124
rect 8067 12121 8079 12155
rect 8021 12115 8079 12121
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 8478 12152 8484 12164
rect 8260 12124 8484 12152
rect 8260 12112 8266 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 10888 12152 10916 12180
rect 10376 12124 10916 12152
rect 10376 12112 10382 12124
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 12618 12152 12624 12164
rect 11112 12124 12624 12152
rect 11112 12112 11118 12124
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 12713 12155 12771 12161
rect 12713 12121 12725 12155
rect 12759 12152 12771 12155
rect 13814 12152 13820 12164
rect 12759 12124 13820 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 15856 12096 15884 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 4338 12044 4344 12096
rect 4396 12044 4402 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5442 12084 5448 12096
rect 4856 12056 5448 12084
rect 4856 12044 4862 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 6730 12084 6736 12096
rect 6512 12056 6736 12084
rect 6512 12044 6518 12056
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 8662 12084 8668 12096
rect 7432 12056 8668 12084
rect 7432 12044 7438 12056
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9214 12084 9220 12096
rect 8812 12056 9220 12084
rect 8812 12044 8818 12056
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 11885 12087 11943 12093
rect 11885 12084 11897 12087
rect 10100 12056 11897 12084
rect 10100 12044 10106 12056
rect 11885 12053 11897 12056
rect 11931 12084 11943 12087
rect 12066 12084 12072 12096
rect 11931 12056 12072 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12253 12087 12311 12093
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 12434 12084 12440 12096
rect 12299 12056 12440 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13170 12084 13176 12096
rect 13127 12056 13176 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13446 12044 13452 12096
rect 13504 12044 13510 12096
rect 15197 12087 15255 12093
rect 15197 12053 15209 12087
rect 15243 12084 15255 12087
rect 15286 12084 15292 12096
rect 15243 12056 15292 12084
rect 15243 12053 15255 12056
rect 15197 12047 15255 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15838 12044 15844 12096
rect 15896 12044 15902 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16224 12084 16252 12183
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16632 12192 16773 12220
rect 16632 12180 16638 12192
rect 16761 12189 16773 12192
rect 16807 12220 16819 12223
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16807 12192 17141 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17236 12220 17264 12328
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 18138 12288 18144 12300
rect 17552 12260 18144 12288
rect 17552 12248 17558 12260
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 17236 12192 17417 12220
rect 17129 12183 17187 12189
rect 17405 12189 17417 12192
rect 17451 12220 17463 12223
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 17451 12192 17693 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 16080 12056 16252 12084
rect 16080 12044 16086 12056
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 17310 12044 17316 12096
rect 17368 12044 17374 12096
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 1104 11994 18860 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 18860 11994
rect 1104 11920 18860 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 6638 11880 6644 11892
rect 2464 11852 6644 11880
rect 2464 11840 2470 11852
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8202 11880 8208 11892
rect 7616 11852 8208 11880
rect 7616 11840 7622 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8662 11880 8668 11892
rect 8343 11852 8668 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9398 11840 9404 11892
rect 9456 11880 9462 11892
rect 9456 11852 10916 11880
rect 9456 11840 9462 11852
rect 3786 11772 3792 11824
rect 3844 11812 3850 11824
rect 4798 11812 4804 11824
rect 3844 11784 4804 11812
rect 3844 11772 3850 11784
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 6788 11784 6837 11812
rect 6788 11772 6794 11784
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 10594 11812 10600 11824
rect 9890 11784 10600 11812
rect 6825 11775 6883 11781
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 10888 11756 10916 11852
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 12216 11852 12265 11880
rect 12216 11840 12222 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 13814 11880 13820 11892
rect 12676 11852 13820 11880
rect 12676 11840 12682 11852
rect 13814 11840 13820 11852
rect 13872 11880 13878 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 13872 11852 14013 11880
rect 13872 11840 13878 11852
rect 14001 11849 14013 11852
rect 14047 11849 14059 11883
rect 14001 11843 14059 11849
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 14148 11852 14657 11880
rect 14148 11840 14154 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 14829 11883 14887 11889
rect 14829 11849 14841 11883
rect 14875 11880 14887 11883
rect 14875 11852 16160 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 11992 11812 12020 11840
rect 13630 11812 13636 11824
rect 11992 11784 13636 11812
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 16025 11815 16083 11821
rect 16025 11781 16037 11815
rect 16071 11781 16083 11815
rect 16132 11812 16160 11852
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 16390 11880 16396 11892
rect 16264 11852 16396 11880
rect 16264 11840 16270 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17310 11812 17316 11824
rect 16132 11784 17316 11812
rect 16025 11775 16083 11781
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2406 11744 2412 11756
rect 2280 11716 2412 11744
rect 2280 11704 2286 11716
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 3050 11744 3056 11756
rect 2639 11716 3056 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6236 11716 6561 11744
rect 6236 11704 6242 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7944 11676 7972 11730
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10502 11744 10508 11756
rect 10459 11716 10508 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 10928 11742 11100 11744
rect 11256 11742 11345 11744
rect 10928 11716 11345 11742
rect 10928 11704 10934 11716
rect 11072 11714 11284 11716
rect 11333 11713 11345 11716
rect 11379 11713 11391 11747
rect 11921 11747 11979 11753
rect 11921 11742 11933 11747
rect 11333 11707 11391 11713
rect 11900 11713 11933 11742
rect 11967 11713 11979 11747
rect 11900 11707 11979 11713
rect 7524 11648 7972 11676
rect 8665 11679 8723 11685
rect 7524 11636 7530 11648
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 8754 11676 8760 11688
rect 8711 11648 8760 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11608 2835 11611
rect 3970 11608 3976 11620
rect 2823 11580 3976 11608
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 6546 11608 6552 11620
rect 5040 11580 6552 11608
rect 5040 11568 5046 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 9968 11608 9996 11704
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 10652 11648 11529 11676
rect 10652 11636 10658 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 11655 11648 11744 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 8220 11580 8524 11608
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 3108 11512 3157 11540
rect 3108 11500 3114 11512
rect 3145 11509 3157 11512
rect 3191 11540 3203 11543
rect 3694 11540 3700 11552
rect 3191 11512 3700 11540
rect 3191 11509 3203 11512
rect 3145 11503 3203 11509
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 8220 11540 8248 11580
rect 4755 11512 8248 11540
rect 8496 11540 8524 11580
rect 9784 11580 9996 11608
rect 10137 11611 10195 11617
rect 9784 11540 9812 11580
rect 10137 11577 10149 11611
rect 10183 11608 10195 11611
rect 11146 11608 11152 11620
rect 10183 11580 11152 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11241 11611 11299 11617
rect 11241 11577 11253 11611
rect 11287 11608 11299 11611
rect 11330 11608 11336 11620
rect 11287 11580 11336 11608
rect 11287 11577 11299 11580
rect 11241 11571 11299 11577
rect 11330 11568 11336 11580
rect 11388 11568 11394 11620
rect 8496 11512 9812 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 9916 11512 10241 11540
rect 9916 11500 9922 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10229 11503 10287 11509
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 10778 11540 10784 11552
rect 10560 11512 10784 11540
rect 10560 11500 10566 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10928 11512 11069 11540
rect 10928 11500 10934 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11716 11540 11744 11648
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 11900 11676 11928 11707
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12216 11716 12265 11744
rect 12216 11704 12222 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 12492 11716 12664 11744
rect 12492 11704 12498 11716
rect 12636 11676 12664 11716
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 13044 11716 15577 11744
rect 13044 11704 13050 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 16040 11744 16068 11775
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 15712 11716 16068 11744
rect 16117 11747 16175 11753
rect 15712 11704 15718 11716
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16206 11744 16212 11756
rect 16163 11716 16212 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16206 11704 16212 11716
rect 16264 11744 16270 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16264 11716 16497 11744
rect 16264 11704 16270 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 13262 11676 13268 11688
rect 11900 11648 12480 11676
rect 12636 11648 13268 11676
rect 11808 11608 11836 11636
rect 12452 11620 12480 11648
rect 13262 11636 13268 11648
rect 13320 11676 13326 11688
rect 14458 11676 14464 11688
rect 13320 11648 14464 11676
rect 13320 11636 13326 11648
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15286 11676 15292 11688
rect 15243 11648 15292 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15841 11679 15899 11685
rect 15841 11645 15853 11679
rect 15887 11676 15899 11679
rect 16022 11676 16028 11688
rect 15887 11648 16028 11676
rect 15887 11645 15899 11648
rect 15841 11639 15899 11645
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 17218 11676 17224 11688
rect 16448 11648 17224 11676
rect 16448 11636 16454 11648
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 11808 11580 11928 11608
rect 11790 11540 11796 11552
rect 11716 11512 11796 11540
rect 11057 11503 11115 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 11900 11540 11928 11580
rect 12434 11568 12440 11620
rect 12492 11568 12498 11620
rect 15562 11568 15568 11620
rect 15620 11568 15626 11620
rect 15654 11568 15660 11620
rect 15712 11568 15718 11620
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 11900 11512 12081 11540
rect 12069 11509 12081 11512
rect 12115 11540 12127 11543
rect 14826 11540 14832 11552
rect 12115 11512 14832 11540
rect 12115 11509 12127 11512
rect 12069 11503 12127 11509
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 1104 11450 18860 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 18860 11450
rect 1104 11376 18860 11398
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6788 11308 6837 11336
rect 6788 11296 6794 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 8018 11336 8024 11348
rect 7147 11308 8024 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10560 11308 10701 11336
rect 10560 11296 10566 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11514 11336 11520 11348
rect 11379 11308 11520 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 4893 11271 4951 11277
rect 4893 11237 4905 11271
rect 4939 11268 4951 11271
rect 5074 11268 5080 11280
rect 4939 11240 5080 11268
rect 4939 11237 4951 11240
rect 4893 11231 4951 11237
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 5258 11228 5264 11280
rect 5316 11268 5322 11280
rect 6549 11271 6607 11277
rect 6549 11268 6561 11271
rect 5316 11240 6561 11268
rect 5316 11228 5322 11240
rect 6549 11237 6561 11240
rect 6595 11237 6607 11271
rect 6549 11231 6607 11237
rect 6638 11228 6644 11280
rect 6696 11228 6702 11280
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 7248 11240 10765 11268
rect 7248 11228 7254 11240
rect 4430 11160 4436 11212
rect 4488 11200 4494 11212
rect 6656 11200 6684 11228
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 4488 11172 6408 11200
rect 6656 11172 9045 11200
rect 4488 11160 4494 11172
rect 6380 11141 6408 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9490 11160 9496 11212
rect 9548 11160 9554 11212
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 10737 11200 10765 11240
rect 11054 11228 11060 11280
rect 11112 11228 11118 11280
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 10560 11172 10640 11200
rect 10737 11172 10885 11200
rect 10560 11160 10566 11172
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6730 11132 6736 11144
rect 6687 11104 6736 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 4724 11064 4752 11095
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7926 11132 7932 11144
rect 7239 11104 7932 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8803 11104 9137 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9125 11101 9137 11104
rect 9171 11132 9183 11135
rect 9214 11132 9220 11144
rect 9171 11104 9220 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 10612 11141 10640 11172
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 11072 11200 11100 11228
rect 10873 11163 10931 11169
rect 10980 11172 11100 11200
rect 10980 11141 11008 11172
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10597 11135 10655 11141
rect 10367 11104 10548 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 9674 11064 9680 11076
rect 4724 11036 9680 11064
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10413 11067 10471 11073
rect 10413 11064 10425 11067
rect 9824 11036 10425 11064
rect 9824 11024 9830 11036
rect 10413 11033 10425 11036
rect 10459 11033 10471 11067
rect 10520 11064 10548 11104
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 10965 11135 11023 11141
rect 10735 11104 10824 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 10796 11064 10824 11104
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 11348 11132 11376 11299
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 12710 11336 12716 11348
rect 12216 11308 12716 11336
rect 12216 11296 12222 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14884 11308 14933 11336
rect 14884 11296 14890 11308
rect 14921 11305 14933 11308
rect 14967 11336 14979 11339
rect 17034 11336 17040 11348
rect 14967 11308 17040 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17586 11336 17592 11348
rect 17359 11308 17592 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 11624 11268 11652 11296
rect 11624 11240 11744 11268
rect 11716 11144 11744 11240
rect 13538 11228 13544 11280
rect 13596 11228 13602 11280
rect 13630 11228 13636 11280
rect 13688 11268 13694 11280
rect 14366 11268 14372 11280
rect 13688 11240 14372 11268
rect 13688 11228 13694 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 17129 11271 17187 11277
rect 17129 11268 17141 11271
rect 15252 11240 17141 11268
rect 15252 11228 15258 11240
rect 17129 11237 17141 11240
rect 17175 11237 17187 11271
rect 17129 11231 17187 11237
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11200 11943 11203
rect 12618 11200 12624 11212
rect 11931 11172 12624 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 13556 11200 13584 11228
rect 13909 11203 13967 11209
rect 13909 11200 13921 11203
rect 13228 11172 13921 11200
rect 13228 11160 13234 11172
rect 13909 11169 13921 11172
rect 13955 11169 13967 11203
rect 13909 11163 13967 11169
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 18138 11200 18144 11212
rect 15887 11172 18144 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 10965 11095 11023 11101
rect 11072 11104 11376 11132
rect 11072 11064 11100 11104
rect 11698 11092 11704 11144
rect 11756 11092 11762 11144
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13596 11104 14105 11132
rect 13596 11092 13602 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14366 11092 14372 11144
rect 14424 11092 14430 11144
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15528 11104 15761 11132
rect 15528 11092 15534 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 16574 11132 16580 11144
rect 15988 11104 16580 11132
rect 15988 11092 15994 11104
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17092 11104 17540 11132
rect 17092 11092 17098 11104
rect 10520 11036 10640 11064
rect 10796 11036 11100 11064
rect 10413 11027 10471 11033
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 7742 10996 7748 11008
rect 6696 10968 7748 10996
rect 6696 10956 6702 10968
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8662 10996 8668 11008
rect 8168 10968 8668 10996
rect 8168 10956 8174 10968
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 10428 10996 10456 11027
rect 10502 10996 10508 11008
rect 10428 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 10612 10996 10640 11036
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 12161 11067 12219 11073
rect 12161 11064 12173 11067
rect 11388 11036 12173 11064
rect 11388 11024 11394 11036
rect 12161 11033 12173 11036
rect 12207 11033 12219 11067
rect 12161 11027 12219 11033
rect 12360 11036 12650 11064
rect 11054 10996 11060 11008
rect 10612 10968 11060 10996
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 11256 10996 11284 11024
rect 12360 11008 12388 11036
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 13872 11036 14197 11064
rect 13872 11024 13878 11036
rect 14185 11033 14197 11036
rect 14231 11033 14243 11067
rect 14185 11027 14243 11033
rect 14553 11067 14611 11073
rect 14553 11033 14565 11067
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 15657 11067 15715 11073
rect 15657 11033 15669 11067
rect 15703 11064 15715 11067
rect 15948 11064 15976 11092
rect 15703 11036 15976 11064
rect 17297 11067 17355 11073
rect 15703 11033 15715 11036
rect 15657 11027 15715 11033
rect 17297 11033 17309 11067
rect 17343 11064 17355 11067
rect 17402 11064 17408 11076
rect 17343 11036 17408 11064
rect 17343 11033 17355 11036
rect 17297 11027 17355 11033
rect 12250 10996 12256 11008
rect 11256 10968 12256 10996
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 14568 10996 14596 11027
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 17512 11073 17540 11104
rect 17497 11067 17555 11073
rect 17497 11033 17509 11067
rect 17543 11033 17555 11067
rect 17497 11027 17555 11033
rect 18506 11024 18512 11076
rect 18564 11024 18570 11076
rect 13136 10968 14596 10996
rect 13136 10956 13142 10968
rect 15470 10956 15476 11008
rect 15528 10996 15534 11008
rect 16022 10996 16028 11008
rect 15528 10968 16028 10996
rect 15528 10956 15534 10968
rect 16022 10956 16028 10968
rect 16080 10996 16086 11008
rect 16209 10999 16267 11005
rect 16209 10996 16221 10999
rect 16080 10968 16221 10996
rect 16080 10956 16086 10968
rect 16209 10965 16221 10968
rect 16255 10965 16267 10999
rect 16209 10959 16267 10965
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17586 10996 17592 11008
rect 17092 10968 17592 10996
rect 17092 10956 17098 10968
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 1104 10906 18860 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 18860 10906
rect 1104 10832 18860 10854
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2372 10764 4568 10792
rect 2372 10752 2378 10764
rect 2498 10616 2504 10668
rect 2556 10656 2562 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2556 10628 2697 10656
rect 2556 10616 2562 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 4540 10656 4568 10764
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 7926 10792 7932 10804
rect 4856 10764 7932 10792
rect 4856 10752 4862 10764
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 8260 10764 9045 10792
rect 8260 10752 8266 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10560 10764 10793 10792
rect 10560 10752 10566 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11885 10795 11943 10801
rect 11388 10764 11744 10792
rect 11388 10752 11394 10764
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 5960 10696 8984 10724
rect 5960 10684 5966 10696
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 2685 10619 2743 10625
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 4080 10588 4108 10642
rect 4540 10628 6377 10656
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 8110 10656 8116 10668
rect 7515 10628 8116 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7190 10588 7196 10600
rect 3007 10560 4016 10588
rect 4080 10560 7196 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3988 10520 4016 10560
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 5442 10520 5448 10532
rect 3988 10492 5448 10520
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 4430 10412 4436 10464
rect 4488 10412 4494 10464
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6420 10424 6561 10452
rect 6420 10412 6426 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 7300 10452 7328 10619
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8772 10588 8800 10619
rect 7984 10560 8800 10588
rect 8956 10588 8984 10696
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 9548 10696 10916 10724
rect 9548 10684 9554 10696
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9122 10656 9128 10668
rect 9079 10628 9128 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9122 10616 9128 10628
rect 9180 10656 9186 10668
rect 9306 10656 9312 10668
rect 9180 10628 9312 10656
rect 9180 10616 9186 10628
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 10888 10656 10916 10696
rect 11514 10684 11520 10736
rect 11572 10684 11578 10736
rect 11716 10733 11744 10764
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 17034 10792 17040 10804
rect 11931 10764 17040 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 11701 10727 11759 10733
rect 11701 10693 11713 10727
rect 11747 10693 11759 10727
rect 12434 10724 12440 10736
rect 11701 10687 11759 10693
rect 12176 10696 12440 10724
rect 12176 10665 12204 10696
rect 12434 10684 12440 10696
rect 12492 10724 12498 10736
rect 15470 10724 15476 10736
rect 12492 10696 15476 10724
rect 12492 10684 12498 10696
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 15930 10684 15936 10736
rect 15988 10724 15994 10736
rect 16206 10724 16212 10736
rect 15988 10696 16212 10724
rect 15988 10684 15994 10696
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 16942 10684 16948 10736
rect 17000 10684 17006 10736
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 10888 10654 11652 10656
rect 11808 10654 11989 10656
rect 10888 10628 11989 10654
rect 11532 10626 11578 10628
rect 11624 10626 11836 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 8956 10560 12081 10588
rect 7984 10548 7990 10560
rect 7653 10523 7711 10529
rect 7653 10489 7665 10523
rect 7699 10520 7711 10523
rect 8570 10520 8576 10532
rect 7699 10492 8576 10520
rect 7699 10489 7711 10492
rect 7653 10483 7711 10489
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7300 10424 7941 10452
rect 6549 10415 6607 10421
rect 7929 10421 7941 10424
rect 7975 10452 7987 10455
rect 8662 10452 8668 10464
rect 7975 10424 8668 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8772 10452 8800 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 8941 10523 8999 10529
rect 8941 10489 8953 10523
rect 8987 10520 8999 10523
rect 11054 10520 11060 10532
rect 8987 10492 11060 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 8772 10424 9321 10452
rect 9309 10421 9321 10424
rect 9355 10452 9367 10455
rect 12176 10452 12204 10619
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 15654 10656 15660 10668
rect 13320 10628 15660 10656
rect 13320 10616 13326 10628
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 16960 10656 16988 10684
rect 17129 10659 17187 10665
rect 17129 10656 17141 10659
rect 16960 10628 17141 10656
rect 17129 10625 17141 10628
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 14734 10588 14740 10600
rect 12308 10560 14740 10588
rect 12308 10548 12314 10560
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 9355 10424 12204 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13136 10424 13921 10452
rect 13136 10412 13142 10424
rect 13909 10421 13921 10424
rect 13955 10452 13967 10455
rect 14458 10452 14464 10464
rect 13955 10424 14464 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17862 10452 17868 10464
rect 17267 10424 17868 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 1104 10362 18860 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 18860 10362
rect 1104 10288 18860 10310
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 14918 10248 14924 10260
rect 4488 10220 14924 10248
rect 4488 10208 4494 10220
rect 14918 10208 14924 10220
rect 14976 10248 14982 10260
rect 15838 10248 15844 10260
rect 14976 10220 15844 10248
rect 14976 10208 14982 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 2314 10140 2320 10192
rect 2372 10180 2378 10192
rect 5994 10180 6000 10192
rect 2372 10152 6000 10180
rect 2372 10140 2378 10152
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 11790 10180 11796 10192
rect 6104 10152 11796 10180
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 3234 9868 3240 9920
rect 3292 9908 3298 9920
rect 3694 9908 3700 9920
rect 3292 9880 3700 9908
rect 3292 9868 3298 9880
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 5718 9868 5724 9920
rect 5776 9868 5782 9920
rect 5920 9908 5948 10007
rect 6104 9985 6132 10152
rect 11790 10140 11796 10152
rect 11848 10180 11854 10192
rect 16206 10180 16212 10192
rect 11848 10152 16212 10180
rect 11848 10140 11854 10152
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 9122 10112 9128 10124
rect 8076 10084 9128 10112
rect 8076 10072 8082 10084
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 10870 10112 10876 10124
rect 10376 10084 10876 10112
rect 10376 10072 10382 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 12342 10112 12348 10124
rect 11020 10084 12348 10112
rect 11020 10072 11026 10084
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18414 10112 18420 10124
rect 18012 10084 18420 10112
rect 18012 10072 18018 10084
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 10594 10044 10600 10056
rect 6227 10016 10600 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6135 9948 6469 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 6457 9939 6515 9945
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 8570 9976 8576 9988
rect 8260 9948 8576 9976
rect 8260 9936 8266 9948
rect 8570 9936 8576 9948
rect 8628 9936 8634 9988
rect 8662 9936 8668 9988
rect 8720 9976 8726 9988
rect 9217 9979 9275 9985
rect 9217 9976 9229 9979
rect 8720 9948 9229 9976
rect 8720 9936 8726 9948
rect 9217 9945 9229 9948
rect 9263 9945 9275 9979
rect 11514 9976 11520 9988
rect 9217 9939 9275 9945
rect 9646 9948 11520 9976
rect 9646 9908 9674 9948
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 5920 9880 9674 9908
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10686 9908 10692 9920
rect 10376 9880 10692 9908
rect 10376 9868 10382 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 12250 9908 12256 9920
rect 10836 9880 12256 9908
rect 10836 9868 10842 9880
rect 12250 9868 12256 9880
rect 12308 9908 12314 9920
rect 15930 9908 15936 9920
rect 12308 9880 15936 9908
rect 12308 9868 12314 9880
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 1104 9818 18860 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 18860 9818
rect 1104 9744 18860 9766
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8478 9704 8484 9716
rect 7064 9676 8484 9704
rect 7064 9664 7070 9676
rect 8478 9664 8484 9676
rect 8536 9704 8542 9716
rect 12618 9704 12624 9716
rect 8536 9676 12624 9704
rect 8536 9664 8542 9676
rect 12618 9664 12624 9676
rect 12676 9704 12682 9716
rect 12897 9707 12955 9713
rect 12897 9704 12909 9707
rect 12676 9676 12909 9704
rect 12676 9664 12682 9676
rect 12897 9673 12909 9676
rect 12943 9673 12955 9707
rect 12897 9667 12955 9673
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 16850 9704 16856 9716
rect 13044 9676 16856 9704
rect 13044 9664 13050 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 4246 9596 4252 9648
rect 4304 9596 4310 9648
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5534 9636 5540 9648
rect 5031 9608 5540 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9398 9596 9404 9648
rect 9456 9596 9462 9648
rect 9766 9596 9772 9648
rect 9824 9636 9830 9648
rect 10778 9636 10784 9648
rect 9824 9608 10784 9636
rect 9824 9596 9830 9608
rect 10778 9596 10784 9608
rect 10836 9636 10842 9648
rect 10836 9608 13216 9636
rect 10836 9596 10842 9608
rect 13188 9580 13216 9608
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 14550 9636 14556 9648
rect 13872 9608 14556 9636
rect 13872 9596 13878 9608
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6420 9540 6960 9568
rect 6420 9528 6426 9540
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 1728 9472 2973 9500
rect 1728 9460 1734 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 6932 9500 6960 9540
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 7742 9568 7748 9580
rect 7699 9540 7748 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6932 9472 7205 9500
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7392 9500 7420 9531
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 10042 9528 10048 9580
rect 10100 9528 10106 9580
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 11900 9540 12357 9568
rect 7558 9500 7564 9512
rect 7392 9472 7564 9500
rect 7193 9463 7251 9469
rect 7558 9460 7564 9472
rect 7616 9500 7622 9512
rect 7616 9472 8156 9500
rect 7616 9460 7622 9472
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 6730 9432 6736 9444
rect 5592 9404 6736 9432
rect 5592 9392 5598 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7285 9435 7343 9441
rect 7285 9401 7297 9435
rect 7331 9401 7343 9435
rect 8128 9432 8156 9472
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9677 9503 9735 9509
rect 9456 9472 9628 9500
rect 9456 9460 9462 9472
rect 8202 9432 8208 9444
rect 8128 9404 8208 9432
rect 7285 9395 7343 9401
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 5960 9336 6837 9364
rect 5960 9324 5966 9336
rect 6825 9333 6837 9336
rect 6871 9364 6883 9367
rect 7006 9364 7012 9376
rect 6871 9336 7012 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7006 9324 7012 9336
rect 7064 9364 7070 9376
rect 7300 9364 7328 9395
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 9600 9432 9628 9472
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 11790 9500 11796 9512
rect 9723 9472 11796 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 11900 9432 11928 9540
rect 12345 9537 12357 9540
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12544 9500 12572 9531
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13078 9568 13084 9580
rect 12676 9540 13084 9568
rect 12676 9528 12682 9540
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 15470 9568 15476 9580
rect 13228 9540 15476 9568
rect 13228 9528 13234 9540
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 16390 9568 16396 9580
rect 15896 9540 16396 9568
rect 15896 9528 15902 9540
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 9600 9404 11928 9432
rect 11992 9472 12572 9500
rect 7064 9336 7328 9364
rect 7561 9367 7619 9373
rect 7064 9324 7070 9336
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 7834 9364 7840 9376
rect 7607 9336 7840 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 10962 9364 10968 9376
rect 8444 9336 10968 9364
rect 8444 9324 8450 9336
rect 10962 9324 10968 9336
rect 11020 9364 11026 9376
rect 11992 9373 12020 9472
rect 12345 9435 12403 9441
rect 12345 9401 12357 9435
rect 12391 9432 12403 9435
rect 16850 9432 16856 9444
rect 12391 9404 16856 9432
rect 12391 9401 12403 9404
rect 12345 9395 12403 9401
rect 16850 9392 16856 9404
rect 16908 9392 16914 9444
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11020 9336 11989 9364
rect 11020 9324 11026 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 11977 9327 12035 9333
rect 1104 9274 18860 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 18860 9274
rect 1104 9200 18860 9222
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 6086 9160 6092 9172
rect 3844 9132 6092 9160
rect 3844 9120 3850 9132
rect 6086 9120 6092 9132
rect 6144 9160 6150 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6144 9132 6285 9160
rect 6144 9120 6150 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 6733 9163 6791 9169
rect 6733 9129 6745 9163
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 5350 9092 5356 9104
rect 2884 9064 5356 9092
rect 2884 8965 2912 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 6748 9092 6776 9123
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 9769 9163 9827 9169
rect 9769 9160 9781 9163
rect 7340 9132 9781 9160
rect 7340 9120 7346 9132
rect 9769 9129 9781 9132
rect 9815 9129 9827 9163
rect 10410 9160 10416 9172
rect 9769 9123 9827 9129
rect 10244 9132 10416 9160
rect 7558 9092 7564 9104
rect 6748 9064 7564 9092
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 8110 9092 8116 9104
rect 7892 9064 8116 9092
rect 7892 9052 7898 9064
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 9033 9095 9091 9101
rect 8251 9064 8892 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 8864 9024 8892 9064
rect 9033 9061 9045 9095
rect 9079 9092 9091 9095
rect 9122 9092 9128 9104
rect 9079 9064 9128 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 10244 9092 10272 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10560 9132 10885 9160
rect 10560 9120 10566 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 10965 9163 11023 9169
rect 10965 9129 10977 9163
rect 11011 9160 11023 9163
rect 11054 9160 11060 9172
rect 11011 9132 11060 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 12032 9132 13737 9160
rect 12032 9120 12038 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 13964 9132 18061 9160
rect 13964 9120 13970 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 10060 9064 10272 9092
rect 10336 9064 10548 9092
rect 9490 9024 9496 9036
rect 4764 8996 7788 9024
rect 4764 8984 4770 8996
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2639 8928 2881 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 4430 8956 4436 8968
rect 3007 8928 4436 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6822 8956 6828 8968
rect 6144 8928 6828 8956
rect 6144 8916 6150 8928
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8956 7619 8959
rect 7650 8956 7656 8968
rect 7607 8928 7656 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 7760 8965 7788 8996
rect 8036 8996 8800 9024
rect 8864 8996 9496 9024
rect 8036 8968 8064 8996
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 8018 8956 8024 8968
rect 7791 8928 8024 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 8662 8956 8668 8968
rect 8343 8928 8668 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 8772 8956 8800 8996
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9674 8984 9680 9036
rect 9732 8984 9738 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10060 9033 10088 9064
rect 9928 9027 9986 9033
rect 9928 9024 9940 9027
rect 9824 8996 9940 9024
rect 9824 8984 9830 8996
rect 9928 8993 9940 8996
rect 9974 8993 9986 9027
rect 9928 8987 9986 8993
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10336 9024 10364 9064
rect 10192 8996 10364 9024
rect 10192 8984 10198 8996
rect 10410 8984 10416 9036
rect 10468 8984 10474 9036
rect 10520 9024 10548 9064
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 11517 9095 11575 9101
rect 11517 9092 11529 9095
rect 10744 9064 11529 9092
rect 10744 9052 10750 9064
rect 10520 8996 10824 9024
rect 10796 8958 10824 8996
rect 11256 8965 11284 9064
rect 11517 9061 11529 9064
rect 11563 9092 11575 9095
rect 11563 9064 12112 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11848 8996 11989 9024
rect 11848 8984 11854 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 12084 9024 12112 9064
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 15562 9092 15568 9104
rect 13504 9064 15568 9092
rect 13504 9052 13510 9064
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 17037 9095 17095 9101
rect 17037 9092 17049 9095
rect 15988 9064 17049 9092
rect 15988 9052 15994 9064
rect 17037 9061 17049 9064
rect 17083 9061 17095 9095
rect 17037 9055 17095 9061
rect 15286 9024 15292 9036
rect 12084 8996 15292 9024
rect 11977 8987 12035 8993
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 10965 8959 11023 8965
rect 10965 8958 10977 8959
rect 8772 8928 10640 8956
rect 10796 8930 10977 8958
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 2464 8860 2697 8888
rect 2464 8848 2470 8860
rect 2685 8857 2697 8860
rect 2731 8857 2743 8891
rect 2685 8851 2743 8857
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 3283 8860 3985 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 3973 8857 3985 8860
rect 4019 8888 4031 8891
rect 4982 8888 4988 8900
rect 4019 8860 4988 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 6730 8888 6736 8900
rect 5592 8860 6736 8888
rect 5592 8848 5598 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7282 8888 7288 8900
rect 7024 8860 7288 8888
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3605 8823 3663 8829
rect 3605 8820 3617 8823
rect 3099 8792 3617 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3605 8789 3617 8792
rect 3651 8820 3663 8823
rect 4062 8820 4068 8832
rect 3651 8792 4068 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 7024 8820 7052 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 7469 8891 7527 8897
rect 7469 8857 7481 8891
rect 7515 8888 7527 8891
rect 9398 8888 9404 8900
rect 7515 8860 9404 8888
rect 7515 8857 7527 8860
rect 7469 8851 7527 8857
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 9784 8860 10517 8888
rect 6420 8792 7052 8820
rect 6420 8780 6426 8792
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7653 8823 7711 8829
rect 7653 8820 7665 8823
rect 7156 8792 7665 8820
rect 7156 8780 7162 8792
rect 7653 8789 7665 8792
rect 7699 8789 7711 8823
rect 7653 8783 7711 8789
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9784 8820 9812 8860
rect 10505 8857 10517 8860
rect 10551 8857 10563 8891
rect 10505 8851 10563 8857
rect 9364 8792 9812 8820
rect 9364 8780 9370 8792
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 10100 8792 10149 8820
rect 10100 8780 10106 8792
rect 10137 8789 10149 8792
rect 10183 8789 10195 8823
rect 10612 8820 10640 8928
rect 10965 8925 10977 8930
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 10686 8848 10692 8900
rect 10744 8848 10750 8900
rect 11164 8888 11192 8919
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14274 8956 14280 8968
rect 13964 8928 14280 8956
rect 13964 8916 13970 8928
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 17052 8956 17080 9055
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17052 8928 17417 8956
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 18064 8956 18092 9123
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18064 8928 18245 8956
rect 17405 8919 17463 8925
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 10796 8860 11192 8888
rect 10796 8820 10824 8860
rect 11422 8848 11428 8900
rect 11480 8888 11486 8900
rect 11882 8888 11888 8900
rect 11480 8860 11888 8888
rect 11480 8848 11486 8860
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 12250 8848 12256 8900
rect 12308 8848 12314 8900
rect 17313 8891 17371 8897
rect 17313 8888 17325 8891
rect 13478 8860 17325 8888
rect 17313 8857 17325 8860
rect 17359 8857 17371 8891
rect 17420 8888 17448 8919
rect 18690 8888 18696 8900
rect 17420 8860 18696 8888
rect 17313 8851 17371 8857
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 10612 8792 10824 8820
rect 10137 8783 10195 8789
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 14274 8820 14280 8832
rect 11204 8792 14280 8820
rect 11204 8780 11210 8792
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 18860 8730
rect 1104 8656 18860 8678
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3786 8616 3792 8628
rect 3467 8588 3792 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 5994 8616 6000 8628
rect 5224 8588 6000 8616
rect 5224 8576 5230 8588
rect 5994 8576 6000 8588
rect 6052 8616 6058 8628
rect 9490 8616 9496 8628
rect 6052 8588 9496 8616
rect 6052 8576 6058 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9582 8576 9588 8628
rect 9640 8576 9646 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 10778 8616 10784 8628
rect 10643 8588 10784 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 11422 8616 11428 8628
rect 11379 8588 11428 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 11422 8576 11428 8588
rect 11480 8616 11486 8628
rect 12529 8619 12587 8625
rect 12529 8616 12541 8619
rect 11480 8588 12541 8616
rect 11480 8576 11486 8588
rect 12529 8585 12541 8588
rect 12575 8616 12587 8619
rect 12986 8616 12992 8628
rect 12575 8588 12992 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 14090 8616 14096 8628
rect 13412 8588 14096 8616
rect 13412 8576 13418 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14182 8576 14188 8628
rect 14240 8576 14246 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14424 8588 18184 8616
rect 14424 8576 14430 8588
rect 3510 8548 3516 8560
rect 3174 8520 3516 8548
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 4172 8548 4200 8576
rect 4893 8551 4951 8557
rect 4893 8548 4905 8551
rect 3804 8520 4905 8548
rect 3804 8489 3832 8520
rect 4893 8517 4905 8520
rect 4939 8517 4951 8551
rect 4893 8511 4951 8517
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 5500 8520 6224 8548
rect 5500 8508 5506 8520
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 3528 8452 3617 8480
rect 3528 8424 3556 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4154 8480 4160 8492
rect 4019 8452 4160 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 1946 8372 1952 8424
rect 2004 8372 2010 8424
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3896 8412 3924 8443
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 6086 8480 6092 8492
rect 5684 8452 6092 8480
rect 5684 8440 5690 8452
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6196 8480 6224 8520
rect 6270 8508 6276 8560
rect 6328 8548 6334 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 6328 8520 6377 8548
rect 6328 8508 6334 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 8021 8551 8079 8557
rect 8021 8517 8033 8551
rect 8067 8517 8079 8551
rect 8021 8511 8079 8517
rect 6196 8452 6776 8480
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 3896 8384 4629 8412
rect 4617 8381 4629 8384
rect 4663 8412 4675 8415
rect 6362 8412 6368 8424
rect 4663 8384 6368 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 6748 8412 6776 8452
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7650 8480 7656 8492
rect 6880 8452 7656 8480
rect 6880 8440 6886 8452
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8036 8424 8064 8511
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 9600 8548 9628 8576
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 8168 8520 9628 8548
rect 9692 8520 10057 8548
rect 8168 8508 8174 8520
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9692 8480 9720 8520
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 10410 8508 10416 8560
rect 10468 8548 10474 8560
rect 10870 8548 10876 8560
rect 10468 8520 10876 8548
rect 10468 8508 10474 8520
rect 10870 8508 10876 8520
rect 10928 8508 10934 8560
rect 12158 8508 12164 8560
rect 12216 8508 12222 8560
rect 12342 8508 12348 8560
rect 12400 8508 12406 8560
rect 13372 8548 13400 8576
rect 18156 8557 18184 8588
rect 12636 8520 13400 8548
rect 18141 8551 18199 8557
rect 9456 8452 9720 8480
rect 10239 8483 10297 8489
rect 9944 8473 10002 8479
rect 9456 8440 9462 8452
rect 9944 8439 9956 8473
rect 9990 8439 10002 8473
rect 10239 8449 10251 8483
rect 10285 8478 10297 8483
rect 12360 8480 12388 8508
rect 10285 8470 10364 8478
rect 10285 8450 10456 8470
rect 10285 8449 10297 8450
rect 10239 8443 10297 8449
rect 10336 8442 10456 8450
rect 9944 8433 10002 8439
rect 6914 8412 6920 8424
rect 6748 8384 6920 8412
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7742 8412 7748 8424
rect 7156 8384 7748 8412
rect 7156 8372 7162 8384
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8018 8372 8024 8424
rect 8076 8372 8082 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9732 8384 9781 8412
rect 9732 8372 9738 8384
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 9959 8356 9987 8433
rect 10428 8356 10456 8442
rect 11716 8452 12388 8480
rect 12437 8483 12495 8489
rect 4249 8347 4307 8353
rect 4249 8313 4261 8347
rect 4295 8344 4307 8347
rect 7834 8344 7840 8356
rect 4295 8316 7840 8344
rect 4295 8313 4307 8316
rect 4249 8307 4307 8313
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 7926 8304 7932 8356
rect 7984 8344 7990 8356
rect 8386 8344 8392 8356
rect 7984 8316 8392 8344
rect 7984 8304 7990 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 9401 8347 9459 8353
rect 9401 8344 9413 8347
rect 9272 8316 9413 8344
rect 9272 8304 9278 8316
rect 9401 8313 9413 8316
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9548 8316 9812 8344
rect 9548 8304 9554 8316
rect 4522 8236 4528 8288
rect 4580 8276 4586 8288
rect 9674 8276 9680 8288
rect 4580 8248 9680 8276
rect 4580 8236 4586 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 9784 8276 9812 8316
rect 9950 8304 9956 8356
rect 10008 8304 10014 8356
rect 10134 8294 10140 8306
rect 10065 8276 10140 8294
rect 9784 8254 10140 8276
rect 10192 8254 10198 8306
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10410 8304 10416 8356
rect 10468 8304 10474 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11716 8344 11744 8452
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12636 8480 12664 8520
rect 18141 8517 18153 8551
rect 18187 8517 18199 8551
rect 18141 8511 18199 8517
rect 12483 8452 12664 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13044 8452 13645 8480
rect 13044 8440 13050 8452
rect 13633 8449 13645 8452
rect 13679 8480 13691 8483
rect 13814 8480 13820 8492
rect 13679 8452 13820 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 11882 8412 11888 8424
rect 11839 8384 11888 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11882 8372 11888 8384
rect 11940 8412 11946 8424
rect 11940 8384 12296 8412
rect 11940 8372 11946 8384
rect 10928 8316 11744 8344
rect 10928 8304 10934 8316
rect 12268 8276 12296 8384
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 14108 8412 14136 8443
rect 14274 8440 14280 8492
rect 14332 8440 14338 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 14792 8452 17417 8480
rect 14792 8440 14798 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 14553 8415 14611 8421
rect 14553 8412 14565 8415
rect 13136 8384 14565 8412
rect 13136 8372 13142 8384
rect 14553 8381 14565 8384
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 12713 8347 12771 8353
rect 12713 8344 12725 8347
rect 12691 8316 12725 8344
rect 12713 8313 12725 8316
rect 12759 8313 12771 8347
rect 12713 8307 12771 8313
rect 12897 8347 12955 8353
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13170 8344 13176 8356
rect 12943 8316 13176 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 12728 8276 12756 8307
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 13504 8316 17509 8344
rect 13504 8304 13510 8316
rect 17497 8313 17509 8316
rect 17543 8313 17555 8347
rect 17497 8307 17555 8313
rect 9784 8248 10180 8254
rect 12268 8248 12756 8276
rect 18417 8279 18475 8285
rect 18417 8245 18429 8279
rect 18463 8276 18475 8279
rect 18506 8276 18512 8288
rect 18463 8248 18512 8276
rect 18463 8245 18475 8248
rect 18417 8239 18475 8245
rect 18506 8236 18512 8248
rect 18564 8236 18570 8288
rect 1104 8186 18860 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 18860 8186
rect 1104 8112 18860 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2179 8044 2789 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2777 8041 2789 8044
rect 2823 8072 2835 8075
rect 3326 8072 3332 8084
rect 2823 8044 3332 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 3927 8044 11192 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4246 7964 4252 8016
rect 4304 7964 4310 8016
rect 6178 7964 6184 8016
rect 6236 7964 6242 8016
rect 6825 8007 6883 8013
rect 6825 7973 6837 8007
rect 6871 8004 6883 8007
rect 11054 8004 11060 8016
rect 6871 7976 11060 8004
rect 6871 7973 6883 7976
rect 6825 7967 6883 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 2976 7908 3832 7936
rect 2976 7880 3004 7908
rect 2958 7868 2964 7880
rect 2746 7840 2964 7868
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 2314 7800 2320 7812
rect 1820 7772 2320 7800
rect 1820 7760 1826 7772
rect 2314 7760 2320 7772
rect 2372 7800 2378 7812
rect 2593 7803 2651 7809
rect 2593 7800 2605 7803
rect 2372 7772 2605 7800
rect 2372 7760 2378 7772
rect 2593 7769 2605 7772
rect 2639 7769 2651 7803
rect 2593 7763 2651 7769
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2746 7732 2774 7840
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3804 7877 3832 7908
rect 4430 7896 4436 7948
rect 4488 7936 4494 7948
rect 6196 7936 6224 7964
rect 8110 7936 8116 7948
rect 4488 7908 8116 7936
rect 4488 7896 4494 7908
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9582 7936 9588 7948
rect 8812 7908 9588 7936
rect 8812 7896 8818 7908
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 10008 7908 10333 7936
rect 10008 7896 10014 7908
rect 10321 7905 10333 7908
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 2809 7803 2867 7809
rect 2809 7769 2821 7803
rect 2855 7800 2867 7803
rect 3418 7800 3424 7812
rect 2855 7772 3424 7800
rect 2855 7769 2867 7772
rect 2809 7763 2867 7769
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 3528 7800 3556 7831
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4304 7840 4813 7868
rect 4304 7828 4310 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 3528 7772 4752 7800
rect 2547 7704 2774 7732
rect 2961 7735 3019 7741
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 4154 7732 4160 7744
rect 3007 7704 4160 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 4724 7741 4752 7772
rect 5074 7760 5080 7812
rect 5132 7760 5138 7812
rect 5534 7760 5540 7812
rect 5592 7760 5598 7812
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 7116 7800 7144 7831
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8294 7868 8300 7880
rect 7708 7840 8300 7868
rect 7708 7828 7714 7840
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10410 7868 10416 7880
rect 10192 7840 10416 7868
rect 10192 7828 10198 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10870 7868 10876 7880
rect 10560 7840 10876 7868
rect 10560 7828 10566 7840
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11164 7854 11192 8044
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 12894 8072 12900 8084
rect 11664 8044 12900 8072
rect 11664 8032 11670 8044
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13722 8072 13728 8084
rect 13587 8044 13728 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 15010 8072 15016 8084
rect 13872 8044 15016 8072
rect 13872 8032 13878 8044
rect 15010 8032 15016 8044
rect 15068 8072 15074 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 15068 8044 17693 8072
rect 15068 8032 15074 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 15286 8004 15292 8016
rect 13188 7976 15292 8004
rect 11790 7896 11796 7948
rect 11848 7936 11854 7948
rect 12529 7939 12587 7945
rect 12529 7936 12541 7939
rect 11848 7908 12541 7936
rect 11848 7896 11854 7908
rect 12529 7905 12541 7908
rect 12575 7905 12587 7939
rect 12529 7899 12587 7905
rect 13188 7877 13216 7976
rect 15286 7964 15292 7976
rect 15344 7964 15350 8016
rect 17696 8004 17724 8035
rect 17696 7976 18092 8004
rect 13264 7908 13492 7936
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 12253 7803 12311 7809
rect 7116 7772 11008 7800
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 5718 7732 5724 7744
rect 4755 7704 5724 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6420 7704 6561 7732
rect 6420 7692 6426 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 6972 7704 7021 7732
rect 6972 7692 6978 7704
rect 7009 7701 7021 7704
rect 7055 7732 7067 7735
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 7055 7704 7389 7732
rect 7055 7701 7067 7704
rect 7009 7695 7067 7701
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 7377 7695 7435 7701
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 8110 7732 8116 7744
rect 7800 7704 8116 7732
rect 7800 7692 7806 7704
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 10778 7692 10784 7744
rect 10836 7692 10842 7744
rect 10980 7732 11008 7772
rect 12253 7769 12265 7803
rect 12299 7800 12311 7803
rect 12710 7800 12716 7812
rect 12299 7772 12716 7800
rect 12299 7769 12311 7772
rect 12253 7763 12311 7769
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 13264 7800 13292 7908
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 12820 7772 13292 7800
rect 11882 7732 11888 7744
rect 10980 7704 11888 7732
rect 11882 7692 11888 7704
rect 11940 7732 11946 7744
rect 12820 7732 12848 7772
rect 11940 7704 12848 7732
rect 11940 7692 11946 7704
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 13372 7732 13400 7831
rect 13464 7800 13492 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 17957 7939 18015 7945
rect 17957 7936 17969 7939
rect 13780 7908 17969 7936
rect 13780 7896 13786 7908
rect 17957 7905 17969 7908
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 13964 7840 14473 7868
rect 13964 7828 13970 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 15010 7868 15016 7880
rect 14691 7840 15016 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 14277 7803 14335 7809
rect 14277 7800 14289 7803
rect 13464 7772 14289 7800
rect 14277 7769 14289 7772
rect 14323 7769 14335 7803
rect 14476 7800 14504 7831
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 18064 7877 18092 7976
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 15804 7840 17877 7868
rect 15804 7828 15810 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 18196 7840 18245 7868
rect 18196 7828 18202 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 14921 7803 14979 7809
rect 14921 7800 14933 7803
rect 14476 7772 14933 7800
rect 14277 7763 14335 7769
rect 14921 7769 14933 7772
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 16942 7800 16948 7812
rect 16724 7772 16948 7800
rect 16724 7760 16730 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 12952 7704 13921 7732
rect 12952 7692 12958 7704
rect 13909 7701 13921 7704
rect 13955 7732 13967 7735
rect 14182 7732 14188 7744
rect 13955 7704 14188 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 14182 7692 14188 7704
rect 14240 7732 14246 7744
rect 14642 7732 14648 7744
rect 14240 7704 14648 7732
rect 14240 7692 14246 7704
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17310 7732 17316 7744
rect 16632 7704 17316 7732
rect 16632 7692 16638 7704
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 18414 7692 18420 7744
rect 18472 7692 18478 7744
rect 1104 7642 18860 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 18860 7642
rect 1104 7568 18860 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2222 7528 2228 7540
rect 1820 7500 2228 7528
rect 1820 7488 1826 7500
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 6822 7528 6828 7540
rect 5092 7500 6828 7528
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 2685 7463 2743 7469
rect 2685 7460 2697 7463
rect 2648 7432 2697 7460
rect 2648 7420 2654 7432
rect 2685 7429 2697 7432
rect 2731 7429 2743 7463
rect 2685 7423 2743 7429
rect 3142 7420 3148 7472
rect 3200 7420 3206 7472
rect 5092 7460 5120 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7524 7500 7849 7528
rect 7524 7488 7530 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 11057 7531 11115 7537
rect 10376 7500 10824 7528
rect 10376 7488 10382 7500
rect 6270 7460 6276 7472
rect 4172 7432 5120 7460
rect 5934 7432 6276 7460
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 1728 7296 2421 7324
rect 1728 7284 1734 7296
rect 2409 7293 2421 7296
rect 2455 7324 2467 7327
rect 3418 7324 3424 7336
rect 2455 7296 3424 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 4172 7333 4200 7432
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 6840 7460 6868 7488
rect 10502 7460 10508 7472
rect 6840 7432 10508 7460
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 7098 7392 7104 7404
rect 5920 7364 7104 7392
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4304 7296 4445 7324
rect 4304 7284 4310 7296
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5350 7324 5356 7336
rect 4755 7296 5356 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 5920 7324 5948 7364
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7892 7364 7941 7392
rect 7892 7352 7898 7364
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 7975 7364 8217 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10413 7395 10471 7401
rect 10413 7392 10425 7395
rect 10376 7364 10425 7392
rect 10376 7352 10382 7364
rect 10413 7361 10425 7364
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 10597 7398 10655 7401
rect 10686 7398 10692 7404
rect 10597 7395 10692 7398
rect 10597 7361 10609 7395
rect 10643 7370 10692 7395
rect 10643 7361 10655 7370
rect 10597 7355 10655 7361
rect 10686 7352 10692 7370
rect 10744 7352 10750 7404
rect 10796 7392 10824 7500
rect 11057 7497 11069 7531
rect 11103 7528 11115 7531
rect 11790 7528 11796 7540
rect 11103 7500 11796 7528
rect 11103 7497 11115 7500
rect 11057 7491 11115 7497
rect 11790 7488 11796 7500
rect 11848 7528 11854 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 11848 7500 12817 7528
rect 11848 7488 11854 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 14918 7488 14924 7540
rect 14976 7488 14982 7540
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 15344 7500 17264 7528
rect 15344 7488 15350 7500
rect 10962 7420 10968 7472
rect 11020 7420 11026 7472
rect 11514 7420 11520 7472
rect 11572 7420 11578 7472
rect 13630 7460 13636 7472
rect 12089 7432 13636 7460
rect 12089 7392 12117 7432
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 15102 7420 15108 7472
rect 15160 7420 15166 7472
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 17129 7463 17187 7469
rect 17129 7460 17141 7463
rect 15436 7432 17141 7460
rect 15436 7420 15442 7432
rect 10796 7364 12117 7392
rect 13354 7352 13360 7404
rect 13412 7392 13418 7404
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 13412 7364 13553 7392
rect 13412 7352 13418 7364
rect 13541 7361 13553 7364
rect 13587 7392 13599 7395
rect 15120 7392 15148 7420
rect 16684 7401 16712 7432
rect 17129 7429 17141 7432
rect 17175 7429 17187 7463
rect 17236 7460 17264 7500
rect 17310 7488 17316 7540
rect 17368 7528 17374 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 17368 7500 17601 7528
rect 17368 7488 17374 7500
rect 17589 7497 17601 7500
rect 17635 7497 17647 7531
rect 17589 7491 17647 7497
rect 17236 7432 17448 7460
rect 17129 7423 17187 7429
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 13587 7364 16405 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 16393 7361 16405 7364
rect 16439 7361 16451 7395
rect 16393 7355 16451 7361
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 16942 7392 16948 7404
rect 16899 7364 16948 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 5776 7296 5948 7324
rect 5776 7284 5782 7296
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 6144 7296 6193 7324
rect 6144 7284 6150 7296
rect 6181 7293 6193 7296
rect 6227 7293 6239 7327
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 6181 7287 6239 7293
rect 6564 7296 10517 7324
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 2498 7188 2504 7200
rect 2372 7160 2504 7188
rect 2372 7148 2378 7160
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 6564 7188 6592 7296
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 13998 7324 14004 7336
rect 10836 7296 14004 7324
rect 10836 7284 10842 7296
rect 13998 7284 14004 7296
rect 14056 7324 14062 7336
rect 15102 7324 15108 7336
rect 14056 7296 15108 7324
rect 14056 7284 14062 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 16408 7324 16436 7355
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 16408 7296 17264 7324
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 12802 7256 12808 7268
rect 7156 7228 12808 7256
rect 7156 7216 7162 7228
rect 12802 7216 12808 7228
rect 12860 7256 12866 7268
rect 13814 7256 13820 7268
rect 12860 7228 13820 7256
rect 12860 7216 12866 7228
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14277 7259 14335 7265
rect 14277 7225 14289 7259
rect 14323 7256 14335 7259
rect 14366 7256 14372 7268
rect 14323 7228 14372 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 14645 7259 14703 7265
rect 14645 7225 14657 7259
rect 14691 7256 14703 7259
rect 14826 7256 14832 7268
rect 14691 7228 14832 7256
rect 14691 7225 14703 7228
rect 14645 7219 14703 7225
rect 14826 7216 14832 7228
rect 14884 7256 14890 7268
rect 15654 7256 15660 7268
rect 14884 7228 15660 7256
rect 14884 7216 14890 7228
rect 15654 7216 15660 7228
rect 15712 7216 15718 7268
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16114 7256 16120 7268
rect 15988 7228 16120 7256
rect 15988 7216 15994 7228
rect 16114 7216 16120 7228
rect 16172 7256 16178 7268
rect 16172 7228 16528 7256
rect 16172 7216 16178 7228
rect 3752 7160 6592 7188
rect 3752 7148 3758 7160
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7466 7188 7472 7200
rect 7064 7160 7472 7188
rect 7064 7148 7070 7160
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 11330 7188 11336 7200
rect 7892 7160 11336 7188
rect 7892 7148 7898 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 13446 7188 13452 7200
rect 12400 7160 13452 7188
rect 12400 7148 12406 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 16298 7188 16304 7200
rect 13688 7160 16304 7188
rect 13688 7148 13694 7160
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16500 7188 16528 7228
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16500 7160 16773 7188
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 17236 7188 17264 7296
rect 17420 7265 17448 7432
rect 17405 7259 17463 7265
rect 17405 7225 17417 7259
rect 17451 7225 17463 7259
rect 17954 7256 17960 7268
rect 17405 7219 17463 7225
rect 17512 7228 17960 7256
rect 17512 7188 17540 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 17236 7160 17540 7188
rect 16761 7151 16819 7157
rect 17586 7148 17592 7200
rect 17644 7148 17650 7200
rect 1104 7098 18860 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 18860 7098
rect 1104 7024 18860 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2682 6984 2688 6996
rect 2372 6956 2688 6984
rect 2372 6944 2378 6956
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 3510 6944 3516 6996
rect 3568 6944 3574 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 7834 6984 7840 6996
rect 5868 6956 7840 6984
rect 5868 6944 5874 6956
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8628 6956 8677 6984
rect 8628 6944 8634 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 9490 6944 9496 6996
rect 9548 6944 9554 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 11609 6987 11667 6993
rect 11609 6984 11621 6987
rect 9640 6956 11621 6984
rect 9640 6944 9646 6956
rect 11609 6953 11621 6956
rect 11655 6953 11667 6987
rect 12158 6984 12164 6996
rect 11609 6947 11667 6953
rect 11808 6956 12164 6984
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 10594 6916 10600 6928
rect 6420 6888 10600 6916
rect 6420 6876 6426 6888
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3568 6820 3985 6848
rect 3568 6808 3574 6820
rect 3973 6817 3985 6820
rect 4019 6848 4031 6851
rect 4246 6848 4252 6860
rect 4019 6820 4252 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 6546 6808 6552 6860
rect 6604 6808 6610 6860
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6932 6789 6960 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10962 6916 10968 6928
rect 10744 6888 10968 6916
rect 10744 6876 10750 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11808 6916 11836 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12526 6984 12532 6996
rect 12483 6956 12532 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12618 6944 12624 6996
rect 12676 6944 12682 6996
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 17129 6987 17187 6993
rect 17129 6984 17141 6987
rect 14056 6956 17141 6984
rect 14056 6944 14062 6956
rect 17129 6953 17141 6956
rect 17175 6984 17187 6987
rect 17586 6984 17592 6996
rect 17175 6956 17592 6984
rect 17175 6953 17187 6956
rect 17129 6947 17187 6953
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 17954 6944 17960 6996
rect 18012 6984 18018 6996
rect 18138 6984 18144 6996
rect 18012 6956 18144 6984
rect 18012 6944 18018 6956
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 13541 6919 13599 6925
rect 13541 6916 13553 6919
rect 11164 6888 11836 6916
rect 11916 6888 13553 6916
rect 9306 6848 9312 6860
rect 7116 6820 9312 6848
rect 7116 6789 7144 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 4028 6684 4261 6712
rect 4028 6672 4034 6684
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 6365 6715 6423 6721
rect 6365 6681 6377 6715
rect 6411 6712 6423 6715
rect 6656 6712 6684 6743
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9416 6780 9444 6811
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9548 6820 10057 6848
rect 9548 6808 9554 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9180 6776 9628 6780
rect 9692 6776 9781 6780
rect 9180 6752 9781 6776
rect 9180 6740 9186 6752
rect 9600 6748 9720 6752
rect 9769 6749 9781 6752
rect 9815 6780 9827 6783
rect 11164 6780 11192 6888
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 9815 6752 11192 6780
rect 11256 6780 11284 6811
rect 11422 6808 11428 6860
rect 11480 6808 11486 6860
rect 11916 6848 11944 6888
rect 13541 6885 13553 6888
rect 13587 6916 13599 6919
rect 14642 6916 14648 6928
rect 13587 6888 14648 6916
rect 13587 6885 13599 6888
rect 13541 6879 13599 6885
rect 14642 6876 14648 6888
rect 14700 6876 14706 6928
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 15378 6916 15384 6928
rect 14976 6888 15384 6916
rect 14976 6876 14982 6888
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 12342 6848 12348 6860
rect 11624 6820 11944 6848
rect 11992 6820 12348 6848
rect 11330 6789 11336 6792
rect 11325 6780 11336 6789
rect 11256 6752 11336 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 11325 6743 11336 6752
rect 11330 6740 11336 6743
rect 11388 6740 11394 6792
rect 11624 6789 11652 6820
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 11757 6783 11815 6789
rect 11757 6749 11769 6783
rect 11803 6780 11815 6783
rect 11803 6749 11836 6780
rect 11757 6743 11836 6749
rect 8938 6712 8944 6724
rect 6411 6684 8944 6712
rect 6411 6681 6423 6684
rect 6365 6675 6423 6681
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 9490 6672 9496 6724
rect 9548 6672 9554 6724
rect 11808 6712 11836 6743
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 11992 6789 12020 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13004 6820 13829 6848
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 13004 6789 13032 6820
rect 13817 6817 13829 6820
rect 13863 6848 13875 6851
rect 13906 6848 13912 6860
rect 13863 6820 13912 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14550 6808 14556 6860
rect 14608 6808 14614 6860
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 14792 6820 15577 6848
rect 14792 6808 14798 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 12989 6783 13047 6789
rect 12989 6782 13001 6783
rect 12912 6780 13001 6782
rect 12492 6754 13001 6780
rect 12492 6752 12940 6754
rect 12492 6740 12498 6752
rect 12989 6749 13001 6754
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 13219 6752 14289 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13832 6724 13860 6752
rect 14277 6749 14289 6752
rect 14323 6780 14335 6783
rect 14826 6780 14832 6792
rect 14323 6752 14832 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 14826 6740 14832 6752
rect 14884 6780 14890 6792
rect 14921 6783 14979 6789
rect 14921 6780 14933 6783
rect 14884 6752 14933 6780
rect 14884 6740 14890 6752
rect 14921 6749 14933 6752
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15010 6740 15016 6792
rect 15068 6740 15074 6792
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 15160 6752 15209 6780
rect 15160 6740 15166 6752
rect 15197 6749 15209 6752
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 15746 6780 15752 6792
rect 15335 6752 15752 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 16022 6740 16028 6792
rect 16080 6740 16086 6792
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 11624 6684 11836 6712
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3050 6644 3056 6656
rect 2556 6616 3056 6644
rect 2556 6604 2562 6616
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 5718 6644 5724 6656
rect 3844 6616 5724 6644
rect 3844 6604 3850 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 7006 6604 7012 6656
rect 7064 6604 7070 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7466 6644 7472 6656
rect 7239 6616 7472 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 8628 6616 9689 6644
rect 8628 6604 8634 6616
rect 9677 6613 9689 6616
rect 9723 6644 9735 6647
rect 10594 6644 10600 6656
rect 9723 6616 10600 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 11330 6644 11336 6656
rect 10919 6616 11336 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 11330 6604 11336 6616
rect 11388 6644 11394 6656
rect 11624 6644 11652 6684
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12308 6684 12940 6712
rect 12308 6672 12314 6684
rect 11388 6616 11652 6644
rect 11388 6604 11394 6616
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 11974 6644 11980 6656
rect 11756 6616 11980 6644
rect 11756 6604 11762 6616
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12216 6616 12449 6644
rect 12216 6604 12222 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 12912 6644 12940 6684
rect 13814 6672 13820 6724
rect 13872 6672 13878 6724
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 14737 6715 14795 6721
rect 14737 6712 14749 6715
rect 14424 6684 14749 6712
rect 14424 6672 14430 6684
rect 14737 6681 14749 6684
rect 14783 6681 14795 6715
rect 14737 6675 14795 6681
rect 15378 6672 15384 6724
rect 15436 6672 15442 6724
rect 16040 6712 16068 6740
rect 17126 6712 17132 6724
rect 15856 6684 17132 6712
rect 13630 6644 13636 6656
rect 12912 6616 13636 6644
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15856 6644 15884 6684
rect 17126 6672 17132 6684
rect 17184 6712 17190 6724
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 17184 6684 17417 6712
rect 17184 6672 17190 6684
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 18506 6712 18512 6724
rect 17405 6675 17463 6681
rect 18064 6684 18512 6712
rect 14700 6616 15884 6644
rect 15933 6647 15991 6653
rect 14700 6604 14706 6616
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16022 6644 16028 6656
rect 15979 6616 16028 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 17420 6644 17448 6675
rect 18064 6656 18092 6684
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 18046 6644 18052 6656
rect 17420 6616 18052 6644
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 18860 6554
rect 1104 6480 18860 6502
rect 3786 6400 3792 6452
rect 3844 6400 3850 6452
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 5626 6440 5632 6452
rect 3927 6412 5632 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 5902 6400 5908 6452
rect 5960 6400 5966 6452
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10226 6440 10232 6452
rect 9907 6412 10232 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11882 6400 11888 6452
rect 11940 6449 11946 6452
rect 11940 6443 11959 6449
rect 11947 6409 11959 6443
rect 11940 6403 11959 6409
rect 11940 6400 11946 6403
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12216 6412 12725 6440
rect 12216 6400 12222 6412
rect 12713 6409 12725 6412
rect 12759 6440 12771 6443
rect 13906 6440 13912 6452
rect 12759 6412 13912 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14148 6412 15148 6440
rect 14148 6400 14154 6412
rect 15120 6384 15148 6412
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 15289 6443 15347 6449
rect 15289 6440 15301 6443
rect 15252 6412 15301 6440
rect 15252 6400 15258 6412
rect 15289 6409 15301 6412
rect 15335 6409 15347 6443
rect 15289 6403 15347 6409
rect 17310 6400 17316 6452
rect 17368 6400 17374 6452
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 3108 6344 6960 6372
rect 3108 6332 3114 6344
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3844 6276 4077 6304
rect 3844 6264 3850 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4430 6304 4436 6316
rect 4295 6276 4436 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4172 6236 4200 6267
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6638 6304 6644 6316
rect 5767 6276 6644 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 4724 6236 4752 6267
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 6932 6304 6960 6344
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 9674 6372 9680 6384
rect 7064 6344 9680 6372
rect 7064 6332 7070 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 11698 6332 11704 6384
rect 11756 6332 11762 6384
rect 13173 6375 13231 6381
rect 13173 6372 13185 6375
rect 11992 6344 13185 6372
rect 11992 6338 12020 6344
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 6932 6276 9781 6304
rect 9769 6273 9781 6276
rect 9815 6304 9827 6307
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9815 6276 10241 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 10229 6273 10241 6276
rect 10275 6304 10287 6307
rect 10778 6304 10784 6316
rect 10275 6276 10784 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11900 6310 12020 6338
rect 13173 6341 13185 6344
rect 13219 6372 13231 6375
rect 13817 6375 13875 6381
rect 13817 6372 13829 6375
rect 13219 6344 13829 6372
rect 13219 6341 13231 6344
rect 13173 6335 13231 6341
rect 13817 6341 13829 6344
rect 13863 6341 13875 6375
rect 13817 6335 13875 6341
rect 14274 6332 14280 6384
rect 14332 6332 14338 6384
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 15473 6375 15531 6381
rect 15473 6372 15485 6375
rect 15160 6344 15485 6372
rect 15160 6332 15166 6344
rect 15473 6341 15485 6344
rect 15519 6341 15531 6375
rect 16114 6372 16120 6384
rect 15473 6335 15531 6341
rect 15672 6344 16120 6372
rect 15672 6316 15700 6344
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 16632 6344 16896 6372
rect 16632 6332 16638 6344
rect 11900 6304 11928 6310
rect 11112 6276 11928 6304
rect 11112 6264 11118 6276
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 12952 6276 13553 6304
rect 12952 6264 12958 6276
rect 13541 6273 13553 6276
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15381 6307 15439 6313
rect 15381 6304 15393 6307
rect 15344 6276 15393 6304
rect 15344 6264 15350 6276
rect 15381 6273 15393 6276
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16666 6264 16672 6316
rect 16724 6264 16730 6316
rect 16868 6313 16896 6344
rect 17126 6332 17132 6384
rect 17184 6372 17190 6384
rect 17184 6344 17264 6372
rect 17184 6332 17190 6344
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17236 6313 17264 6344
rect 17402 6332 17408 6384
rect 17460 6372 17466 6384
rect 17460 6344 18000 6372
rect 17460 6332 17466 6344
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 17972 6313 18000 6344
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 17552 6276 17693 6304
rect 17552 6264 17558 6276
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18138 6264 18144 6316
rect 18196 6264 18202 6316
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18325 6307 18383 6313
rect 18325 6304 18337 6307
rect 18288 6276 18337 6304
rect 18288 6264 18294 6276
rect 18325 6273 18337 6276
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 4798 6236 4804 6248
rect 4172 6208 4292 6236
rect 4724 6208 4804 6236
rect 4264 6180 4292 6208
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6236 4951 6239
rect 8846 6236 8852 6248
rect 4939 6208 8852 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 10502 6236 10508 6248
rect 8996 6208 10508 6236
rect 8996 6196 9002 6208
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 11698 6236 11704 6248
rect 10652 6208 11704 6236
rect 10652 6196 10658 6208
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 13814 6236 13820 6248
rect 11900 6208 13820 6236
rect 4246 6128 4252 6180
rect 4304 6128 4310 6180
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 4479 6140 5549 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 5537 6137 5549 6140
rect 5583 6168 5595 6171
rect 7466 6168 7472 6180
rect 5583 6140 7472 6168
rect 5583 6137 5595 6140
rect 5537 6131 5595 6137
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4580 6072 5181 6100
rect 4580 6060 4586 6072
rect 5169 6069 5181 6072
rect 5215 6100 5227 6103
rect 5994 6100 6000 6112
rect 5215 6072 6000 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 11330 6100 11336 6112
rect 6880 6072 11336 6100
rect 6880 6060 6886 6072
rect 11330 6060 11336 6072
rect 11388 6100 11394 6112
rect 11900 6109 11928 6208
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 16684 6236 16712 6264
rect 17405 6239 17463 6245
rect 16684 6208 17264 6236
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 12345 6171 12403 6177
rect 12345 6168 12357 6171
rect 12216 6140 12357 6168
rect 12216 6128 12222 6140
rect 12345 6137 12357 6140
rect 12391 6168 12403 6171
rect 12618 6168 12624 6180
rect 12391 6140 12624 6168
rect 12391 6137 12403 6140
rect 12345 6131 12403 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13078 6168 13084 6180
rect 12768 6140 13084 6168
rect 12768 6128 12774 6140
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6168 15899 6171
rect 16666 6168 16672 6180
rect 15887 6140 16672 6168
rect 15887 6137 15899 6140
rect 15841 6131 15899 6137
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 16850 6128 16856 6180
rect 16908 6128 16914 6180
rect 17236 6168 17264 6208
rect 17405 6205 17417 6239
rect 17451 6236 17463 6239
rect 17770 6236 17776 6248
rect 17451 6208 17776 6236
rect 17451 6205 17463 6208
rect 17405 6199 17463 6205
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 18141 6171 18199 6177
rect 18141 6168 18153 6171
rect 17236 6140 18153 6168
rect 18141 6137 18153 6140
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11388 6072 11897 6100
rect 11388 6060 11394 6072
rect 11885 6069 11897 6072
rect 11931 6069 11943 6103
rect 11885 6063 11943 6069
rect 12066 6060 12072 6112
rect 12124 6060 12130 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12526 6100 12532 6112
rect 12308 6072 12532 6100
rect 12308 6060 12314 6072
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12636 6100 12664 6128
rect 13814 6100 13820 6112
rect 12636 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 16114 6060 16120 6112
rect 16172 6060 16178 6112
rect 1104 6010 18860 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 18860 6010
rect 1104 5936 18860 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3234 5896 3240 5908
rect 2823 5868 3240 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3694 5896 3700 5908
rect 3559 5868 3700 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3528 5828 3556 5859
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4614 5896 4620 5908
rect 4571 5868 4620 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 4724 5868 5825 5896
rect 2148 5800 3556 5828
rect 2148 5769 2176 5800
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 4724 5828 4752 5868
rect 5813 5865 5825 5868
rect 5859 5896 5871 5899
rect 7374 5896 7380 5908
rect 5859 5868 7380 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7432 5868 8033 5896
rect 7432 5856 7438 5868
rect 8021 5865 8033 5868
rect 8067 5896 8079 5899
rect 9766 5896 9772 5908
rect 8067 5868 9772 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 10836 5868 11253 5896
rect 10836 5856 10842 5868
rect 11241 5865 11253 5868
rect 11287 5865 11299 5899
rect 11241 5859 11299 5865
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12584 5868 12817 5896
rect 12584 5856 12590 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 13078 5856 13084 5908
rect 13136 5856 13142 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5865 13323 5899
rect 13265 5859 13323 5865
rect 4488 5800 4752 5828
rect 4488 5788 4494 5800
rect 4798 5788 4804 5840
rect 4856 5788 4862 5840
rect 5077 5831 5135 5837
rect 5077 5797 5089 5831
rect 5123 5828 5135 5831
rect 5442 5828 5448 5840
rect 5123 5800 5448 5828
rect 5123 5797 5135 5800
rect 5077 5791 5135 5797
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 5776 5800 9444 5828
rect 5776 5788 5782 5800
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 3142 5760 3148 5772
rect 2133 5723 2191 5729
rect 2608 5732 3148 5760
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2608 5701 2636 5732
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 4816 5760 4844 5788
rect 4816 5732 5488 5760
rect 5460 5704 5488 5732
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 4062 5692 4068 5704
rect 2823 5664 4068 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 9416 5692 9444 5800
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 13280 5828 13308 5859
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 15197 5899 15255 5905
rect 15197 5896 15209 5899
rect 15160 5868 15209 5896
rect 15160 5856 15166 5868
rect 15197 5865 15209 5868
rect 15243 5865 15255 5899
rect 15197 5859 15255 5865
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 15565 5899 15623 5905
rect 15565 5896 15577 5899
rect 15344 5868 15577 5896
rect 15344 5856 15350 5868
rect 15565 5865 15577 5868
rect 15611 5865 15623 5899
rect 17218 5896 17224 5908
rect 15565 5859 15623 5865
rect 16316 5868 17224 5896
rect 10928 5800 13308 5828
rect 10928 5788 10934 5800
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 13630 5828 13636 5840
rect 13412 5800 13636 5828
rect 13412 5788 13418 5800
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 16316 5837 16344 5868
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17402 5856 17408 5908
rect 17460 5856 17466 5908
rect 17865 5899 17923 5905
rect 17865 5865 17877 5899
rect 17911 5896 17923 5899
rect 18230 5896 18236 5908
rect 17911 5868 18236 5896
rect 17911 5865 17923 5868
rect 17865 5859 17923 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 14384 5800 16313 5828
rect 14384 5772 14412 5800
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 12618 5760 12624 5772
rect 9548 5732 12624 5760
rect 9548 5720 9554 5732
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 14366 5760 14372 5772
rect 12820 5732 14372 5760
rect 9766 5692 9772 5704
rect 9416 5664 9772 5692
rect 9766 5652 9772 5664
rect 9824 5692 9830 5704
rect 10042 5692 10048 5704
rect 9824 5664 10048 5692
rect 9824 5652 9830 5664
rect 10042 5652 10048 5664
rect 10100 5692 10106 5704
rect 12820 5692 12848 5732
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5760 14979 5763
rect 15654 5760 15660 5772
rect 14967 5732 15660 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 16574 5720 16580 5772
rect 16632 5720 16638 5772
rect 10100 5664 12848 5692
rect 10100 5652 10106 5664
rect 12894 5652 12900 5704
rect 12952 5692 12958 5704
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 12952 5664 13553 5692
rect 12952 5652 12958 5664
rect 13541 5661 13553 5664
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 16592 5692 16620 5720
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 13964 5664 16681 5692
rect 13964 5652 13970 5664
rect 16669 5661 16681 5664
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 17552 5664 18245 5692
rect 17552 5652 17558 5664
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 6362 5624 6368 5636
rect 4939 5596 6368 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 9582 5624 9588 5636
rect 8352 5596 9588 5624
rect 8352 5584 8358 5596
rect 9582 5584 9588 5596
rect 9640 5624 9646 5636
rect 9953 5627 10011 5633
rect 9953 5624 9965 5627
rect 9640 5596 9965 5624
rect 9640 5584 9646 5596
rect 9953 5593 9965 5596
rect 9999 5593 10011 5627
rect 9953 5587 10011 5593
rect 10594 5584 10600 5636
rect 10652 5584 10658 5636
rect 10778 5584 10784 5636
rect 10836 5633 10842 5636
rect 10836 5627 10855 5633
rect 10843 5593 10855 5627
rect 12802 5624 12808 5636
rect 10836 5587 10855 5593
rect 10888 5596 12808 5624
rect 10836 5584 10842 5587
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 4062 5556 4068 5568
rect 2547 5528 4068 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4430 5556 4436 5568
rect 4304 5528 4436 5556
rect 4304 5516 4310 5528
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 10888 5556 10916 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13262 5633 13268 5636
rect 13249 5627 13268 5633
rect 13249 5624 13261 5627
rect 13136 5596 13261 5624
rect 13136 5584 13142 5596
rect 13249 5593 13261 5596
rect 13249 5587 13268 5593
rect 13262 5584 13268 5587
rect 13320 5584 13326 5636
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 13412 5596 13461 5624
rect 13412 5584 13418 5596
rect 13449 5593 13461 5596
rect 13495 5593 13507 5627
rect 13449 5587 13507 5593
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5624 13783 5627
rect 13814 5624 13820 5636
rect 13771 5596 13820 5624
rect 13771 5593 13783 5596
rect 13725 5587 13783 5593
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 15746 5584 15752 5636
rect 15804 5624 15810 5636
rect 17037 5627 17095 5633
rect 17037 5624 17049 5627
rect 15804 5596 17049 5624
rect 15804 5584 15810 5596
rect 17037 5593 17049 5596
rect 17083 5624 17095 5627
rect 17126 5624 17132 5636
rect 17083 5596 17132 5624
rect 17083 5593 17095 5596
rect 17037 5587 17095 5593
rect 17126 5584 17132 5596
rect 17184 5624 17190 5636
rect 17770 5624 17776 5636
rect 17184 5596 17776 5624
rect 17184 5584 17190 5596
rect 17770 5584 17776 5596
rect 17828 5584 17834 5636
rect 10560 5528 10916 5556
rect 10560 5516 10566 5528
rect 10962 5516 10968 5568
rect 11020 5516 11026 5568
rect 18414 5516 18420 5568
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 2685 5355 2743 5361
rect 2685 5352 2697 5355
rect 1636 5324 2697 5352
rect 1636 5312 1642 5324
rect 2685 5321 2697 5324
rect 2731 5321 2743 5355
rect 2685 5315 2743 5321
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7432 5324 7481 5352
rect 7432 5312 7438 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 9306 5352 9312 5364
rect 7469 5315 7527 5321
rect 8128 5324 9312 5352
rect 2406 5244 2412 5296
rect 2464 5244 2470 5296
rect 4430 5244 4436 5296
rect 4488 5284 4494 5296
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 4488 5256 7297 5284
rect 4488 5244 4494 5256
rect 7285 5253 7297 5256
rect 7331 5284 7343 5287
rect 8128 5284 8156 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 9640 5324 10333 5352
rect 9640 5312 9646 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 13078 5352 13084 5364
rect 10836 5324 13084 5352
rect 10836 5312 10842 5324
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 13633 5355 13691 5361
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 13814 5352 13820 5364
rect 13679 5324 13820 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13906 5312 13912 5364
rect 13964 5312 13970 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16669 5355 16727 5361
rect 15896 5324 16436 5352
rect 15896 5312 15902 5324
rect 7331 5256 8156 5284
rect 7331 5253 7343 5256
rect 7285 5247 7343 5253
rect 2498 5176 2504 5228
rect 2556 5216 2562 5228
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2556 5188 2605 5216
rect 2556 5176 2562 5188
rect 2593 5185 2605 5188
rect 2639 5216 2651 5219
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 2639 5188 3065 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 3053 5185 3065 5188
rect 3099 5216 3111 5219
rect 5810 5216 5816 5228
rect 3099 5188 5816 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 7392 5225 7420 5256
rect 8202 5244 8208 5296
rect 8260 5284 8266 5296
rect 8297 5287 8355 5293
rect 8297 5284 8309 5287
rect 8260 5256 8309 5284
rect 8260 5244 8266 5256
rect 8297 5253 8309 5256
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 9030 5244 9036 5296
rect 9088 5244 9094 5296
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10137 5287 10195 5293
rect 10137 5284 10149 5287
rect 10008 5256 10149 5284
rect 10008 5244 10014 5256
rect 10137 5253 10149 5256
rect 10183 5284 10195 5287
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10183 5256 10701 5284
rect 10183 5253 10195 5256
rect 10137 5247 10195 5253
rect 10689 5253 10701 5256
rect 10735 5284 10747 5287
rect 11606 5284 11612 5296
rect 10735 5256 11612 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7423 5188 7457 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7616 5188 7665 5216
rect 7616 5176 7622 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 4246 5148 4252 5160
rect 1912 5120 4252 5148
rect 1912 5108 1918 5120
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 7668 5148 7696 5179
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10318 5216 10324 5228
rect 10091 5188 10324 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 15930 5216 15936 5228
rect 10459 5188 15936 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 11330 5148 11336 5160
rect 7668 5120 11336 5148
rect 11330 5108 11336 5120
rect 11388 5148 11394 5160
rect 16408 5148 16436 5324
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16758 5352 16764 5364
rect 16715 5324 16764 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5321 17095 5355
rect 17037 5315 17095 5321
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 17052 5284 17080 5315
rect 17218 5312 17224 5364
rect 17276 5312 17282 5364
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 18141 5355 18199 5361
rect 18141 5352 18153 5355
rect 18104 5324 18153 5352
rect 18104 5312 18110 5324
rect 18141 5321 18153 5324
rect 18187 5321 18199 5355
rect 18141 5315 18199 5321
rect 16540 5256 17080 5284
rect 16540 5244 16546 5256
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 17494 5216 17500 5228
rect 16632 5188 17500 5216
rect 16632 5176 16638 5188
rect 17494 5176 17500 5188
rect 17552 5216 17558 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17552 5188 17785 5216
rect 17552 5176 17558 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 11388 5120 16865 5148
rect 11388 5108 11394 5120
rect 16853 5117 16865 5120
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 16942 5108 16948 5160
rect 17000 5108 17006 5160
rect 17126 5108 17132 5160
rect 17184 5148 17190 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 17184 5120 17325 5148
rect 17184 5108 17190 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 9364 5052 10088 5080
rect 9364 5040 9370 5052
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 6822 5012 6828 5024
rect 2363 4984 6828 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 9950 5012 9956 5024
rect 7883 4984 9956 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10060 5012 10088 5052
rect 10134 5040 10140 5092
rect 10192 5040 10198 5092
rect 10318 5040 10324 5092
rect 10376 5080 10382 5092
rect 10376 5052 13308 5080
rect 10376 5040 10382 5052
rect 13280 5024 13308 5052
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 17144 5080 17172 5108
rect 16632 5052 17172 5080
rect 16632 5040 16638 5052
rect 13078 5012 13084 5024
rect 10060 4984 13084 5012
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 16114 5012 16120 5024
rect 15528 4984 16120 5012
rect 15528 4972 15534 4984
rect 16114 4972 16120 4984
rect 16172 5012 16178 5024
rect 16942 5012 16948 5024
rect 16172 4984 16948 5012
rect 16172 4972 16178 4984
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 1104 4922 18860 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 18860 4922
rect 1104 4848 18860 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 1820 4780 3985 4808
rect 1820 4768 1826 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 3973 4771 4031 4777
rect 4338 4768 4344 4820
rect 4396 4768 4402 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 6822 4808 6828 4820
rect 5040 4780 6828 4808
rect 5040 4768 5046 4780
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 7193 4811 7251 4817
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 7282 4808 7288 4820
rect 7239 4780 7288 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 7024 4740 7052 4771
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7616 4780 8125 4808
rect 7616 4768 7622 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 10318 4808 10324 4820
rect 8536 4780 10324 4808
rect 8536 4768 8542 4780
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 10652 4780 12541 4808
rect 10652 4768 10658 4780
rect 12529 4777 12541 4780
rect 12575 4777 12587 4811
rect 12529 4771 12587 4777
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 15194 4808 15200 4820
rect 13136 4780 15200 4808
rect 13136 4768 13142 4780
rect 15194 4768 15200 4780
rect 15252 4808 15258 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15252 4780 16129 4808
rect 15252 4768 15258 4780
rect 16117 4777 16129 4780
rect 16163 4808 16175 4811
rect 16482 4808 16488 4820
rect 16163 4780 16488 4808
rect 16163 4777 16175 4780
rect 16117 4771 16175 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16574 4768 16580 4820
rect 16632 4768 16638 4820
rect 16850 4768 16856 4820
rect 16908 4808 16914 4820
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 16908 4780 17049 4808
rect 16908 4768 16914 4780
rect 17037 4777 17049 4780
rect 17083 4777 17095 4811
rect 17037 4771 17095 4777
rect 17221 4811 17279 4817
rect 17221 4777 17233 4811
rect 17267 4808 17279 4811
rect 18322 4808 18328 4820
rect 17267 4780 18328 4808
rect 17267 4777 17279 4780
rect 17221 4771 17279 4777
rect 7374 4740 7380 4752
rect 7024 4712 7380 4740
rect 7374 4700 7380 4712
rect 7432 4740 7438 4752
rect 8570 4740 8576 4752
rect 7432 4712 8576 4740
rect 7432 4700 7438 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 10229 4743 10287 4749
rect 10229 4709 10241 4743
rect 10275 4740 10287 4743
rect 10410 4740 10416 4752
rect 10275 4712 10416 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 10686 4700 10692 4752
rect 10744 4740 10750 4752
rect 10781 4743 10839 4749
rect 10781 4740 10793 4743
rect 10744 4712 10793 4740
rect 10744 4700 10750 4712
rect 10781 4709 10793 4712
rect 10827 4709 10839 4743
rect 10781 4703 10839 4709
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 12161 4743 12219 4749
rect 12161 4740 12173 4743
rect 11204 4712 12173 4740
rect 11204 4700 11210 4712
rect 12161 4709 12173 4712
rect 12207 4740 12219 4743
rect 14645 4743 14703 4749
rect 12207 4712 12434 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6917 4675 6975 4681
rect 6917 4672 6929 4675
rect 6144 4644 6929 4672
rect 6144 4632 6150 4644
rect 6917 4641 6929 4644
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8352 4644 10272 4672
rect 8352 4632 8358 4644
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 4338 4604 4344 4616
rect 3835 4576 4344 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6236 4576 6745 4604
rect 6236 4564 6242 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6880 4576 7021 4604
rect 6880 4564 6886 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7466 4604 7472 4616
rect 7055 4576 7472 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8680 4576 9076 4604
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 8680 4536 8708 4576
rect 5868 4508 8708 4536
rect 8757 4539 8815 4545
rect 5868 4496 5874 4508
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8803 4508 8953 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 9048 4536 9076 4576
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9640 4576 9812 4604
rect 9640 4564 9646 4576
rect 9677 4539 9735 4545
rect 9677 4536 9689 4539
rect 9048 4508 9689 4536
rect 8941 4499 8999 4505
rect 9677 4505 9689 4508
rect 9723 4505 9735 4539
rect 9784 4536 9812 4576
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10244 4613 10272 4644
rect 10612 4644 12296 4672
rect 10612 4613 10640 4644
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 11146 4536 11152 4548
rect 9784 4508 11152 4536
rect 9677 4499 9735 4505
rect 8956 4468 8984 4499
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 10870 4468 10876 4480
rect 8956 4440 10876 4468
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 12268 4468 12296 4644
rect 12406 4604 12434 4712
rect 14645 4709 14657 4743
rect 14691 4740 14703 4743
rect 15102 4740 15108 4752
rect 14691 4712 15108 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 15286 4700 15292 4752
rect 15344 4740 15350 4752
rect 15565 4743 15623 4749
rect 15565 4740 15577 4743
rect 15344 4712 15577 4740
rect 15344 4700 15350 4712
rect 15565 4709 15577 4712
rect 15611 4709 15623 4743
rect 15565 4703 15623 4709
rect 13446 4672 13452 4684
rect 13188 4644 13452 4672
rect 13188 4613 13216 4644
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12406 4576 12725 4604
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12943 4576 13185 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13262 4564 13268 4616
rect 13320 4604 13326 4616
rect 17052 4604 17080 4771
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18141 4743 18199 4749
rect 18141 4709 18153 4743
rect 18187 4740 18199 4743
rect 18690 4740 18696 4752
rect 18187 4712 18696 4740
rect 18187 4709 18199 4712
rect 18141 4703 18199 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 13320 4576 15424 4604
rect 17052 4576 17417 4604
rect 13320 4564 13326 4576
rect 14918 4496 14924 4548
rect 14976 4496 14982 4548
rect 15102 4496 15108 4548
rect 15160 4496 15166 4548
rect 15286 4496 15292 4548
rect 15344 4496 15350 4548
rect 15396 4536 15424 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 17773 4539 17831 4545
rect 17773 4536 17785 4539
rect 15396 4508 17785 4536
rect 17773 4505 17785 4508
rect 17819 4536 17831 4539
rect 18138 4536 18144 4548
rect 17819 4508 18144 4536
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 15010 4468 15016 4480
rect 12268 4440 15016 4468
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 18414 4428 18420 4480
rect 18472 4428 18478 4480
rect 1104 4378 18860 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 18860 4378
rect 1104 4304 18860 4326
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 3878 4264 3884 4276
rect 2087 4236 3884 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 6362 4264 6368 4276
rect 4120 4236 6368 4264
rect 4120 4224 4126 4236
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7374 4224 7380 4276
rect 7432 4224 7438 4276
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8478 4264 8484 4276
rect 8435 4236 8484 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 8662 4273 8668 4276
rect 8649 4267 8668 4273
rect 8649 4233 8661 4267
rect 8649 4227 8668 4233
rect 8662 4224 8668 4227
rect 8720 4224 8726 4276
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11112 4236 11897 4264
rect 11112 4224 11118 4236
rect 11885 4233 11897 4236
rect 11931 4233 11943 4267
rect 11885 4227 11943 4233
rect 12621 4267 12679 4273
rect 12621 4233 12633 4267
rect 12667 4264 12679 4267
rect 13998 4264 14004 4276
rect 12667 4236 14004 4264
rect 12667 4233 12679 4236
rect 12621 4227 12679 4233
rect 2498 4196 2504 4208
rect 1872 4168 2504 4196
rect 1872 4140 1900 4168
rect 2498 4156 2504 4168
rect 2556 4156 2562 4208
rect 4246 4156 4252 4208
rect 4304 4156 4310 4208
rect 8294 4196 8300 4208
rect 5474 4168 8300 4196
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 8496 4196 8524 4224
rect 8849 4199 8907 4205
rect 8849 4196 8861 4199
rect 8496 4168 8861 4196
rect 8849 4165 8861 4168
rect 8895 4196 8907 4199
rect 8938 4196 8944 4208
rect 8895 4168 8944 4196
rect 8895 4165 8907 4168
rect 8849 4159 8907 4165
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 9030 4156 9036 4208
rect 9088 4196 9094 4208
rect 9674 4196 9680 4208
rect 9088 4168 9680 4196
rect 9088 4156 9094 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 10042 4156 10048 4208
rect 10100 4156 10106 4208
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 11204 4168 11529 4196
rect 11204 4156 11210 4168
rect 11517 4165 11529 4168
rect 11563 4165 11575 4199
rect 11517 4159 11575 4165
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11733 4199 11791 4205
rect 11733 4196 11745 4199
rect 11664 4168 11745 4196
rect 11664 4156 11670 4168
rect 11733 4165 11745 4168
rect 11779 4196 11791 4199
rect 12636 4196 12664 4227
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 17497 4267 17555 4273
rect 17497 4264 17509 4267
rect 15620 4236 17509 4264
rect 15620 4224 15626 4236
rect 17497 4233 17509 4236
rect 17543 4264 17555 4267
rect 18023 4267 18081 4273
rect 18023 4264 18035 4267
rect 17543 4236 18035 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 18023 4233 18035 4236
rect 18069 4233 18081 4267
rect 18023 4227 18081 4233
rect 11779 4168 12664 4196
rect 13357 4199 13415 4205
rect 11779 4165 11791 4168
rect 11733 4159 11791 4165
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13722 4196 13728 4208
rect 13403 4168 13728 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 18138 4156 18144 4208
rect 18196 4196 18202 4208
rect 18233 4199 18291 4205
rect 18233 4196 18245 4199
rect 18196 4168 18245 4196
rect 18196 4156 18202 4168
rect 18233 4165 18245 4168
rect 18279 4165 18291 4199
rect 18233 4159 18291 4165
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2271 4100 2774 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 1762 3884 1768 3936
rect 1820 3884 1826 3936
rect 2424 3924 2452 4023
rect 2746 3992 2774 4100
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6788 4100 8524 4128
rect 6788 4088 6794 4100
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3970 4060 3976 4072
rect 3568 4032 3976 4060
rect 3568 4020 3574 4032
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4614 4060 4620 4072
rect 4080 4032 4620 4060
rect 4080 3992 4108 4032
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 2746 3964 4108 3992
rect 6549 3995 6607 4001
rect 6549 3961 6561 3995
rect 6595 3992 6607 3995
rect 8202 3992 8208 4004
rect 6595 3964 8208 3992
rect 6595 3961 6607 3964
rect 6549 3955 6607 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 8496 4001 8524 4100
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 18325 4131 18383 4137
rect 13219 4100 13768 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3961 8539 3995
rect 8481 3955 8539 3961
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2424 3896 2697 3924
rect 2685 3893 2697 3896
rect 2731 3924 2743 3927
rect 6822 3924 6828 3936
rect 2731 3896 6828 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8168 3896 8677 3924
rect 8168 3884 8174 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 9324 3924 9352 4023
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11333 4063 11391 4069
rect 11333 4060 11345 4063
rect 11296 4032 11345 4060
rect 11296 4020 11302 4032
rect 11333 4029 11345 4032
rect 11379 4060 11391 4063
rect 11790 4060 11796 4072
rect 11379 4032 11796 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 13740 4069 13768 4100
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 18690 4128 18696 4140
rect 18371 4100 18696 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 14826 4060 14832 4072
rect 13771 4032 14832 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 16724 3964 18092 3992
rect 16724 3952 16730 3964
rect 9582 3924 9588 3936
rect 9324 3896 9588 3924
rect 8665 3887 8723 3893
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 10226 3924 10232 3936
rect 9640 3896 10232 3924
rect 9640 3884 9646 3896
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11747 3896 12173 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 12161 3893 12173 3896
rect 12207 3924 12219 3927
rect 13538 3924 13544 3936
rect 12207 3896 13544 3924
rect 12207 3893 12219 3896
rect 12161 3887 12219 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 17862 3884 17868 3936
rect 17920 3884 17926 3936
rect 18064 3933 18092 3964
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18196 3896 18429 3924
rect 18196 3884 18202 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 1104 3834 18860 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 18860 3834
rect 1104 3760 18860 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1912 3692 1961 3720
rect 1912 3680 1918 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 2958 3680 2964 3732
rect 3016 3680 3022 3732
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 5534 3720 5540 3732
rect 3283 3692 5540 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 9125 3723 9183 3729
rect 6512 3692 8064 3720
rect 6512 3680 6518 3692
rect 8036 3652 8064 3692
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 12066 3720 12072 3732
rect 9171 3692 12072 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 16448 3692 17601 3720
rect 16448 3680 16454 3692
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 9490 3652 9496 3664
rect 8036 3624 9496 3652
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 11330 3612 11336 3664
rect 11388 3612 11394 3664
rect 12345 3655 12403 3661
rect 12345 3621 12357 3655
rect 12391 3652 12403 3655
rect 13814 3652 13820 3664
rect 12391 3624 13820 3652
rect 12391 3621 12403 3624
rect 12345 3615 12403 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 4028 3556 6745 3584
rect 4028 3544 4034 3556
rect 6733 3553 6745 3556
rect 6779 3584 6791 3587
rect 8018 3584 8024 3596
rect 6779 3556 8024 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9582 3584 9588 3596
rect 9272 3556 9588 3584
rect 9272 3544 9278 3556
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9858 3544 9864 3596
rect 9916 3544 9922 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10008 3556 12204 3584
rect 10008 3544 10014 3556
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 3016 3488 3157 3516
rect 3016 3476 3022 3488
rect 3145 3485 3157 3488
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 9490 3516 9496 3528
rect 8803 3488 9496 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11164 3488 11621 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 5316 3420 7021 3448
rect 5316 3408 5322 3420
rect 7009 3417 7021 3420
rect 7055 3417 7067 3451
rect 8662 3448 8668 3460
rect 8234 3420 8668 3448
rect 7009 3411 7067 3417
rect 8662 3408 8668 3420
rect 8720 3408 8726 3460
rect 8938 3408 8944 3460
rect 8996 3408 9002 3460
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9141 3451 9199 3457
rect 9141 3448 9153 3451
rect 9088 3420 9153 3448
rect 9088 3408 9094 3420
rect 9141 3417 9153 3420
rect 9187 3417 9199 3451
rect 9950 3448 9956 3460
rect 9141 3411 9199 3417
rect 9232 3420 9956 3448
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 9232 3380 9260 3420
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 4212 3352 9260 3380
rect 4212 3340 4218 3352
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 11164 3380 11192 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11698 3476 11704 3528
rect 11756 3476 11762 3528
rect 11790 3476 11796 3528
rect 11848 3476 11854 3528
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 12176 3525 12204 3556
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3485 12219 3519
rect 17604 3516 17632 3683
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17604 3488 17785 3516
rect 12161 3479 12219 3485
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18782 3516 18788 3528
rect 18279 3488 18788 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 17310 3448 17316 3460
rect 12084 3420 17316 3448
rect 11514 3380 11520 3392
rect 9456 3352 11520 3380
rect 9456 3340 9462 3352
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 12084 3389 12112 3420
rect 17310 3408 17316 3420
rect 17368 3408 17374 3460
rect 12069 3383 12127 3389
rect 12069 3349 12081 3383
rect 12115 3349 12127 3383
rect 12069 3343 12127 3349
rect 12158 3340 12164 3392
rect 12216 3380 12222 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 12216 3352 12633 3380
rect 12216 3340 12222 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 12986 3340 12992 3392
rect 13044 3340 13050 3392
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 16264 3352 17877 3380
rect 16264 3340 16270 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 18414 3340 18420 3392
rect 18472 3340 18478 3392
rect 1104 3290 18860 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 18860 3290
rect 1104 3216 18860 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 10042 3176 10048 3188
rect 1820 3148 10048 3176
rect 1820 3136 1826 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 10870 3176 10876 3188
rect 10367 3148 10876 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 11756 3148 12541 3176
rect 11756 3136 11762 3148
rect 12529 3145 12541 3148
rect 12575 3176 12587 3179
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 12575 3148 13185 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14424 3148 14565 3176
rect 14424 3136 14430 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 15102 3176 15108 3188
rect 15059 3148 15108 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 15102 3136 15108 3148
rect 15160 3176 15166 3188
rect 15746 3176 15752 3188
rect 15160 3148 15752 3176
rect 15160 3136 15166 3148
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3108 8907 3111
rect 8938 3108 8944 3120
rect 8895 3080 8944 3108
rect 8895 3077 8907 3080
rect 8849 3071 8907 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 10560 3080 10609 3108
rect 10560 3068 10566 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 10597 3071 10655 3077
rect 11514 3068 11520 3120
rect 11572 3068 11578 3120
rect 11808 3080 12020 3108
rect 11808 3052 11836 3080
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 8720 3012 10824 3040
rect 8720 3000 8726 3012
rect 10796 2972 10824 3012
rect 10870 3000 10876 3052
rect 10928 3000 10934 3052
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 11882 3000 11888 3052
rect 11940 3000 11946 3052
rect 11992 3040 12020 3080
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 12434 3108 12440 3120
rect 12124 3080 12440 3108
rect 12124 3068 12130 3080
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 11992 3012 12817 3040
rect 12805 3009 12817 3012
rect 12851 3040 12863 3043
rect 12986 3040 12992 3052
rect 12851 3012 12992 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 10796 2944 12434 2972
rect 11241 2907 11299 2913
rect 11241 2904 11253 2907
rect 6104 2876 11253 2904
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 6104 2845 6132 2876
rect 11241 2873 11253 2876
rect 11287 2904 11299 2907
rect 11882 2904 11888 2916
rect 11287 2876 11888 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 11882 2864 11888 2876
rect 11940 2904 11946 2916
rect 12158 2904 12164 2916
rect 11940 2876 12164 2904
rect 11940 2864 11946 2876
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12406 2904 12434 2944
rect 17402 2904 17408 2916
rect 12406 2876 17408 2904
rect 17402 2864 17408 2876
rect 17460 2864 17466 2916
rect 6089 2839 6147 2845
rect 6089 2836 6101 2839
rect 5592 2808 6101 2836
rect 5592 2796 5598 2808
rect 6089 2805 6101 2808
rect 6135 2805 6147 2839
rect 6089 2799 6147 2805
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 8386 2836 8392 2848
rect 6880 2808 8392 2836
rect 6880 2796 6886 2808
rect 8386 2796 8392 2808
rect 8444 2836 8450 2848
rect 12069 2839 12127 2845
rect 12069 2836 12081 2839
rect 8444 2808 12081 2836
rect 8444 2796 8450 2808
rect 12069 2805 12081 2808
rect 12115 2805 12127 2839
rect 12069 2799 12127 2805
rect 1104 2746 18860 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 18860 2746
rect 1104 2672 18860 2694
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2632 6699 2635
rect 11241 2635 11299 2641
rect 6687 2604 11192 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 6656 2564 6684 2595
rect 6104 2536 6684 2564
rect 11164 2564 11192 2604
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11422 2632 11428 2644
rect 11287 2604 11428 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 14737 2635 14795 2641
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 15194 2632 15200 2644
rect 14783 2604 15200 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 11698 2564 11704 2576
rect 11164 2536 11704 2564
rect 5534 2388 5540 2440
rect 5592 2388 5598 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6104 2428 6132 2536
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 14918 2524 14924 2576
rect 14976 2524 14982 2576
rect 9490 2456 9496 2508
rect 9548 2456 9554 2508
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 15381 2499 15439 2505
rect 15381 2496 15393 2499
rect 14415 2468 15393 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 15381 2465 15393 2468
rect 15427 2496 15439 2499
rect 16114 2496 16120 2508
rect 15427 2468 16120 2496
rect 15427 2465 15439 2468
rect 15381 2459 15439 2465
rect 16114 2456 16120 2468
rect 16172 2456 16178 2508
rect 5859 2400 6132 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 3660 2332 9137 2360
rect 3660 2320 3666 2332
rect 9125 2329 9137 2332
rect 9171 2360 9183 2363
rect 9769 2363 9827 2369
rect 9769 2360 9781 2363
rect 9171 2332 9781 2360
rect 9171 2329 9183 2332
rect 9125 2323 9183 2329
rect 9769 2329 9781 2332
rect 9815 2329 9827 2363
rect 13170 2360 13176 2372
rect 10994 2332 13176 2360
rect 9769 2323 9827 2329
rect 13170 2320 13176 2332
rect 13228 2320 13234 2372
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 15212 2360 15240 2391
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18598 2428 18604 2440
rect 18279 2400 18604 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 14424 2332 15240 2360
rect 14424 2320 14430 2332
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 5675 2264 7021 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 7009 2261 7021 2264
rect 7055 2292 7067 2295
rect 11790 2292 11796 2304
rect 7055 2264 11796 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 18414 2252 18420 2304
rect 18472 2252 18478 2304
rect 1104 2202 18860 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 7288 17552 7340 17604
rect 15660 17552 15712 17604
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 9772 17280 9824 17332
rect 10508 17280 10560 17332
rect 18512 17323 18564 17332
rect 18512 17289 18521 17323
rect 18521 17289 18555 17323
rect 18555 17289 18564 17323
rect 18512 17280 18564 17289
rect 8484 17255 8536 17264
rect 8484 17221 8493 17255
rect 8493 17221 8527 17255
rect 8527 17221 8536 17255
rect 8484 17212 8536 17221
rect 9680 17212 9732 17264
rect 13452 17212 13504 17264
rect 3424 17008 3476 17060
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7748 17187 7800 17196
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 10600 17144 10652 17196
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 14372 17144 14424 17196
rect 15660 17255 15712 17264
rect 15660 17221 15669 17255
rect 15669 17221 15703 17255
rect 15703 17221 15712 17255
rect 15660 17212 15712 17221
rect 7288 17076 7340 17085
rect 3148 16940 3200 16992
rect 4252 16983 4304 16992
rect 4252 16949 4261 16983
rect 4261 16949 4295 16983
rect 4295 16949 4304 16983
rect 4252 16940 4304 16949
rect 11612 17076 11664 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 10876 17008 10928 17060
rect 11704 16940 11756 16992
rect 13268 16940 13320 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14648 16983 14700 16992
rect 14648 16949 14657 16983
rect 14657 16949 14691 16983
rect 14691 16949 14700 16983
rect 14648 16940 14700 16949
rect 16764 16940 16816 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 1768 16736 1820 16788
rect 4252 16736 4304 16788
rect 14004 16736 14056 16788
rect 3148 16668 3200 16720
rect 3792 16668 3844 16720
rect 1676 16532 1728 16584
rect 3792 16532 3844 16584
rect 5080 16600 5132 16652
rect 7472 16668 7524 16720
rect 14648 16668 14700 16720
rect 4344 16464 4396 16516
rect 5264 16532 5316 16584
rect 11704 16600 11756 16652
rect 4252 16396 4304 16448
rect 4988 16439 5040 16448
rect 4988 16405 4997 16439
rect 4997 16405 5031 16439
rect 5031 16405 5040 16439
rect 4988 16396 5040 16405
rect 5632 16396 5684 16448
rect 9220 16532 9272 16584
rect 6092 16464 6144 16516
rect 7748 16464 7800 16516
rect 8300 16464 8352 16516
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 11796 16396 11848 16448
rect 13176 16600 13228 16652
rect 14188 16643 14240 16652
rect 14188 16609 14197 16643
rect 14197 16609 14231 16643
rect 14231 16609 14240 16643
rect 14188 16600 14240 16609
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 12532 16507 12584 16516
rect 12532 16473 12541 16507
rect 12541 16473 12575 16507
rect 12575 16473 12584 16507
rect 12532 16464 12584 16473
rect 15660 16532 15712 16584
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14832 16464 14884 16516
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 8208 16192 8260 16244
rect 10692 16192 10744 16244
rect 5816 16124 5868 16176
rect 5908 16167 5960 16176
rect 5908 16133 5917 16167
rect 5917 16133 5951 16167
rect 5951 16133 5960 16167
rect 5908 16124 5960 16133
rect 6000 16124 6052 16176
rect 8116 16124 8168 16176
rect 15200 16124 15252 16176
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 14832 16056 14884 16108
rect 15476 16056 15528 16108
rect 6184 16031 6236 16040
rect 6184 15997 6193 16031
rect 6193 15997 6227 16031
rect 6227 15997 6236 16031
rect 6184 15988 6236 15997
rect 6368 15988 6420 16040
rect 11244 15988 11296 16040
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 3792 15852 3844 15904
rect 5816 15852 5868 15904
rect 12624 15852 12676 15904
rect 17408 15988 17460 16040
rect 14464 15852 14516 15904
rect 14740 15852 14792 15904
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 16304 15852 16356 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 6368 15648 6420 15700
rect 3884 15580 3936 15632
rect 8208 15648 8260 15700
rect 8760 15648 8812 15700
rect 2504 15512 2556 15564
rect 6184 15512 6236 15564
rect 6368 15512 6420 15564
rect 6644 15512 6696 15564
rect 7288 15512 7340 15564
rect 8024 15512 8076 15564
rect 1584 15444 1636 15496
rect 4436 15444 4488 15496
rect 4620 15444 4672 15496
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 9588 15580 9640 15632
rect 10416 15580 10468 15632
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 13176 15648 13228 15700
rect 15844 15648 15896 15700
rect 12624 15580 12676 15632
rect 13360 15580 13412 15632
rect 16580 15580 16632 15632
rect 2136 15419 2188 15428
rect 2136 15385 2145 15419
rect 2145 15385 2179 15419
rect 2179 15385 2188 15419
rect 2136 15376 2188 15385
rect 2412 15308 2464 15360
rect 4068 15308 4120 15360
rect 4712 15419 4764 15428
rect 4712 15385 4721 15419
rect 4721 15385 4755 15419
rect 4755 15385 4764 15419
rect 4712 15376 4764 15385
rect 4896 15419 4948 15428
rect 4896 15385 4905 15419
rect 4905 15385 4939 15419
rect 4939 15385 4948 15419
rect 4896 15376 4948 15385
rect 6000 15376 6052 15428
rect 7840 15419 7892 15428
rect 7840 15385 7867 15419
rect 7867 15385 7892 15419
rect 7840 15376 7892 15385
rect 8024 15419 8076 15428
rect 8024 15385 8033 15419
rect 8033 15385 8067 15419
rect 8067 15385 8076 15419
rect 8024 15376 8076 15385
rect 10324 15444 10376 15496
rect 11060 15512 11112 15564
rect 9588 15376 9640 15428
rect 11244 15444 11296 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 15292 15512 15344 15564
rect 14464 15444 14516 15496
rect 13636 15376 13688 15428
rect 15660 15376 15712 15428
rect 5264 15308 5316 15360
rect 8484 15308 8536 15360
rect 9404 15308 9456 15360
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 15016 15308 15068 15360
rect 15568 15308 15620 15360
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 13728 15104 13780 15156
rect 14004 15147 14056 15156
rect 14004 15113 14031 15147
rect 14031 15113 14056 15147
rect 14004 15104 14056 15113
rect 15200 15147 15252 15156
rect 15200 15113 15209 15147
rect 15209 15113 15243 15147
rect 15243 15113 15252 15147
rect 15200 15104 15252 15113
rect 1584 15079 1636 15088
rect 1584 15045 1593 15079
rect 1593 15045 1627 15079
rect 1627 15045 1636 15079
rect 1584 15036 1636 15045
rect 6092 15036 6144 15088
rect 6460 15036 6512 15088
rect 9312 15036 9364 15088
rect 9496 15079 9548 15088
rect 9496 15045 9523 15079
rect 9523 15045 9548 15079
rect 9496 15036 9548 15045
rect 10140 15036 10192 15088
rect 14188 15079 14240 15088
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 14832 15036 14884 15088
rect 15568 15036 15620 15088
rect 5724 14968 5776 15020
rect 2320 14764 2372 14816
rect 10324 14900 10376 14952
rect 10600 14900 10652 14952
rect 10876 14900 10928 14952
rect 4160 14832 4212 14884
rect 5724 14832 5776 14884
rect 6368 14832 6420 14884
rect 6184 14764 6236 14816
rect 8392 14764 8444 14816
rect 9128 14764 9180 14816
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 10692 14764 10744 14816
rect 12348 14764 12400 14816
rect 13912 14764 13964 14816
rect 16488 14900 16540 14952
rect 16028 14832 16080 14884
rect 14832 14764 14884 14816
rect 18604 14764 18656 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 3516 14560 3568 14612
rect 4344 14560 4396 14612
rect 6460 14560 6512 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 7380 14560 7432 14612
rect 7748 14560 7800 14612
rect 5724 14492 5776 14544
rect 6000 14492 6052 14544
rect 9404 14560 9456 14612
rect 13360 14560 13412 14612
rect 1676 14356 1728 14408
rect 5080 14424 5132 14476
rect 5172 14424 5224 14476
rect 7472 14424 7524 14476
rect 8116 14424 8168 14476
rect 11980 14424 12032 14476
rect 12072 14424 12124 14476
rect 2320 14356 2372 14408
rect 2412 14356 2464 14408
rect 3792 14356 3844 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5080 14288 5132 14340
rect 2320 14220 2372 14272
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 12440 14356 12492 14408
rect 13544 14424 13596 14476
rect 14372 14424 14424 14476
rect 15752 14424 15804 14476
rect 17316 14492 17368 14544
rect 17500 14424 17552 14476
rect 15108 14356 15160 14408
rect 18880 14356 18932 14408
rect 7748 14220 7800 14272
rect 8116 14331 8168 14340
rect 8116 14297 8125 14331
rect 8125 14297 8159 14331
rect 8159 14297 8168 14331
rect 8116 14288 8168 14297
rect 11244 14288 11296 14340
rect 15292 14288 15344 14340
rect 16856 14288 16908 14340
rect 11336 14220 11388 14272
rect 16212 14220 16264 14272
rect 16396 14220 16448 14272
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 4068 13948 4120 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 4896 14016 4948 14068
rect 4988 14016 5040 14068
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 5172 13948 5224 14000
rect 5540 13948 5592 14000
rect 6000 13948 6052 14000
rect 6460 13948 6512 14000
rect 7288 14016 7340 14068
rect 8668 14016 8720 14068
rect 11980 14016 12032 14068
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 16212 14016 16264 14068
rect 2412 13812 2464 13864
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 6184 13880 6236 13932
rect 9404 13948 9456 14000
rect 11428 13948 11480 14000
rect 12348 13948 12400 14000
rect 13268 13948 13320 14000
rect 14096 13991 14148 14000
rect 14096 13957 14105 13991
rect 14105 13957 14139 13991
rect 14139 13957 14148 13991
rect 14096 13948 14148 13957
rect 15752 13948 15804 14000
rect 13544 13880 13596 13932
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 15200 13880 15252 13932
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 17960 14016 18012 14068
rect 5080 13812 5132 13864
rect 5172 13812 5224 13864
rect 7472 13812 7524 13864
rect 8944 13812 8996 13864
rect 10416 13812 10468 13864
rect 4896 13676 4948 13728
rect 6000 13676 6052 13728
rect 6460 13676 6512 13728
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 6644 13676 6696 13728
rect 9680 13676 9732 13728
rect 10140 13676 10192 13728
rect 12716 13744 12768 13796
rect 12808 13744 12860 13796
rect 13268 13744 13320 13796
rect 15660 13812 15712 13864
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 17316 13812 17368 13864
rect 18144 13855 18196 13864
rect 18144 13821 18153 13855
rect 18153 13821 18187 13855
rect 18187 13821 18196 13855
rect 18144 13812 18196 13821
rect 12348 13676 12400 13728
rect 12900 13676 12952 13728
rect 16304 13676 16356 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 4436 13472 4488 13524
rect 4988 13472 5040 13524
rect 5448 13472 5500 13524
rect 4896 13336 4948 13388
rect 6184 13336 6236 13388
rect 3884 13311 3936 13320
rect 3884 13277 3893 13311
rect 3893 13277 3927 13311
rect 3927 13277 3936 13311
rect 3884 13268 3936 13277
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 6828 13404 6880 13456
rect 12900 13472 12952 13524
rect 8116 13336 8168 13388
rect 10324 13336 10376 13388
rect 5172 13200 5224 13252
rect 6460 13200 6512 13252
rect 7380 13268 7432 13320
rect 9956 13268 10008 13320
rect 8208 13200 8260 13252
rect 9036 13200 9088 13252
rect 16120 13472 16172 13524
rect 17408 13472 17460 13524
rect 17592 13472 17644 13524
rect 17868 13472 17920 13524
rect 17960 13472 18012 13524
rect 18144 13472 18196 13524
rect 13728 13336 13780 13388
rect 14648 13336 14700 13388
rect 15108 13336 15160 13388
rect 18144 13336 18196 13388
rect 13820 13268 13872 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 3608 13132 3660 13184
rect 6644 13132 6696 13184
rect 6736 13132 6788 13184
rect 6920 13132 6972 13184
rect 7564 13132 7616 13184
rect 12808 13132 12860 13184
rect 13636 13200 13688 13252
rect 16580 13200 16632 13252
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 6828 12928 6880 12980
rect 3700 12903 3752 12912
rect 3700 12869 3709 12903
rect 3709 12869 3743 12903
rect 3743 12869 3752 12903
rect 3700 12860 3752 12869
rect 6184 12860 6236 12912
rect 7748 12860 7800 12912
rect 2964 12792 3016 12844
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 3792 12792 3844 12844
rect 1768 12724 1820 12776
rect 10048 12928 10100 12980
rect 8576 12860 8628 12912
rect 10968 12860 11020 12912
rect 11520 12928 11572 12980
rect 3056 12699 3108 12708
rect 3056 12665 3065 12699
rect 3065 12665 3099 12699
rect 3099 12665 3108 12699
rect 3056 12656 3108 12665
rect 4068 12656 4120 12708
rect 6000 12656 6052 12708
rect 7748 12656 7800 12708
rect 5540 12588 5592 12640
rect 6368 12588 6420 12640
rect 7564 12588 7616 12640
rect 8852 12724 8904 12776
rect 10324 12724 10376 12776
rect 10784 12792 10836 12844
rect 15568 12860 15620 12912
rect 15936 12860 15988 12912
rect 16304 12860 16356 12912
rect 16580 12860 16632 12912
rect 11704 12792 11756 12844
rect 12440 12792 12492 12844
rect 12900 12792 12952 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 15292 12792 15344 12844
rect 18052 12792 18104 12844
rect 9312 12656 9364 12708
rect 9588 12631 9640 12640
rect 9588 12597 9597 12631
rect 9597 12597 9631 12631
rect 9631 12597 9640 12631
rect 9588 12588 9640 12597
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11796 12631 11848 12640
rect 11152 12588 11204 12597
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 12256 12588 12308 12640
rect 13912 12699 13964 12708
rect 13912 12665 13921 12699
rect 13921 12665 13955 12699
rect 13955 12665 13964 12699
rect 13912 12656 13964 12665
rect 14648 12724 14700 12776
rect 15476 12724 15528 12776
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 16672 12656 16724 12708
rect 17592 12588 17644 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 2228 12384 2280 12436
rect 3516 12384 3568 12436
rect 4436 12316 4488 12368
rect 6000 12384 6052 12436
rect 7564 12384 7616 12436
rect 8024 12384 8076 12436
rect 9220 12384 9272 12436
rect 9864 12384 9916 12436
rect 10324 12384 10376 12436
rect 11704 12384 11756 12436
rect 11888 12384 11940 12436
rect 14372 12384 14424 12436
rect 16856 12384 16908 12436
rect 16948 12384 17000 12436
rect 17500 12384 17552 12436
rect 17592 12384 17644 12436
rect 18236 12384 18288 12436
rect 3516 12248 3568 12300
rect 3884 12180 3936 12232
rect 4344 12180 4396 12232
rect 6644 12316 6696 12368
rect 8300 12316 8352 12368
rect 12164 12316 12216 12368
rect 12624 12316 12676 12368
rect 6184 12248 6236 12300
rect 7472 12248 7524 12300
rect 12256 12248 12308 12300
rect 2412 12087 2464 12096
rect 3792 12155 3844 12164
rect 3792 12121 3801 12155
rect 3801 12121 3835 12155
rect 3835 12121 3844 12155
rect 3792 12112 3844 12121
rect 10600 12180 10652 12232
rect 10876 12180 10928 12232
rect 11428 12180 11480 12232
rect 11704 12180 11756 12232
rect 12808 12180 12860 12232
rect 13268 12180 13320 12232
rect 13452 12180 13504 12232
rect 14372 12180 14424 12232
rect 14556 12180 14608 12232
rect 2412 12053 2437 12087
rect 2437 12053 2464 12087
rect 2412 12044 2464 12053
rect 3976 12044 4028 12096
rect 6920 12112 6972 12164
rect 8208 12112 8260 12164
rect 8484 12112 8536 12164
rect 10324 12112 10376 12164
rect 11060 12112 11112 12164
rect 12624 12112 12676 12164
rect 13820 12112 13872 12164
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 5448 12044 5500 12096
rect 6460 12044 6512 12096
rect 6736 12044 6788 12096
rect 7380 12044 7432 12096
rect 8668 12044 8720 12096
rect 8760 12044 8812 12096
rect 9220 12044 9272 12096
rect 10048 12044 10100 12096
rect 12072 12044 12124 12096
rect 12440 12044 12492 12096
rect 13176 12044 13228 12096
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 15292 12044 15344 12096
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 16028 12044 16080 12096
rect 16580 12180 16632 12232
rect 17500 12248 17552 12300
rect 18144 12248 18196 12300
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 2412 11840 2464 11892
rect 6644 11840 6696 11892
rect 7564 11840 7616 11892
rect 8208 11840 8260 11892
rect 8668 11840 8720 11892
rect 9404 11840 9456 11892
rect 3792 11772 3844 11824
rect 4804 11772 4856 11824
rect 6736 11772 6788 11824
rect 10600 11772 10652 11824
rect 11980 11840 12032 11892
rect 12164 11840 12216 11892
rect 12624 11840 12676 11892
rect 13820 11840 13872 11892
rect 14096 11840 14148 11892
rect 13636 11772 13688 11824
rect 16212 11840 16264 11892
rect 16396 11840 16448 11892
rect 2228 11704 2280 11756
rect 2412 11704 2464 11756
rect 3056 11704 3108 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 6184 11704 6236 11756
rect 7472 11636 7524 11688
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 9956 11704 10008 11756
rect 10508 11704 10560 11756
rect 10876 11704 10928 11756
rect 8760 11636 8812 11688
rect 3976 11568 4028 11620
rect 4988 11568 5040 11620
rect 6552 11568 6604 11620
rect 10600 11636 10652 11688
rect 3056 11500 3108 11552
rect 3700 11500 3752 11552
rect 11152 11568 11204 11620
rect 11336 11568 11388 11620
rect 9864 11500 9916 11552
rect 10508 11500 10560 11552
rect 10784 11500 10836 11552
rect 10876 11500 10928 11552
rect 11796 11636 11848 11688
rect 12164 11704 12216 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 12992 11704 13044 11756
rect 15660 11704 15712 11756
rect 17316 11772 17368 11824
rect 16212 11704 16264 11756
rect 13268 11636 13320 11688
rect 14464 11636 14516 11688
rect 15292 11636 15344 11688
rect 16028 11636 16080 11688
rect 16396 11636 16448 11688
rect 17224 11636 17276 11688
rect 11796 11500 11848 11552
rect 12440 11568 12492 11620
rect 15568 11611 15620 11620
rect 15568 11577 15577 11611
rect 15577 11577 15611 11611
rect 15611 11577 15620 11611
rect 15568 11568 15620 11577
rect 15660 11611 15712 11620
rect 15660 11577 15669 11611
rect 15669 11577 15703 11611
rect 15703 11577 15712 11611
rect 15660 11568 15712 11577
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 6736 11296 6788 11348
rect 8024 11296 8076 11348
rect 10508 11296 10560 11348
rect 5080 11228 5132 11280
rect 5264 11228 5316 11280
rect 6644 11228 6696 11280
rect 7196 11228 7248 11280
rect 4436 11160 4488 11212
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 10508 11160 10560 11212
rect 11060 11228 11112 11280
rect 6736 11092 6788 11144
rect 7932 11092 7984 11144
rect 9220 11092 9272 11144
rect 9680 11024 9732 11076
rect 9772 11024 9824 11076
rect 11520 11296 11572 11348
rect 11612 11296 11664 11348
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 12164 11296 12216 11348
rect 12716 11296 12768 11348
rect 14832 11296 14884 11348
rect 17040 11296 17092 11348
rect 17592 11296 17644 11348
rect 13544 11228 13596 11280
rect 13636 11228 13688 11280
rect 14372 11228 14424 11280
rect 15200 11228 15252 11280
rect 12624 11160 12676 11212
rect 13176 11160 13228 11212
rect 18144 11160 18196 11212
rect 11704 11092 11756 11144
rect 13544 11092 13596 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15476 11092 15528 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16580 11092 16632 11144
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 6644 10956 6696 11008
rect 7748 10956 7800 11008
rect 8116 10956 8168 11008
rect 8668 10956 8720 11008
rect 10508 10956 10560 11008
rect 11244 11024 11296 11076
rect 11336 11024 11388 11076
rect 11060 10956 11112 11008
rect 13820 11024 13872 11076
rect 12256 10956 12308 11008
rect 12348 10956 12400 11008
rect 13084 10956 13136 11008
rect 17408 11024 17460 11076
rect 18512 11067 18564 11076
rect 18512 11033 18521 11067
rect 18521 11033 18555 11067
rect 18555 11033 18564 11067
rect 18512 11024 18564 11033
rect 15476 10956 15528 11008
rect 16028 10956 16080 11008
rect 17040 10956 17092 11008
rect 17592 10956 17644 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 2320 10752 2372 10804
rect 2504 10616 2556 10668
rect 4804 10752 4856 10804
rect 7932 10752 7984 10804
rect 8208 10752 8260 10804
rect 10508 10752 10560 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 5908 10684 5960 10736
rect 7196 10548 7248 10600
rect 5448 10480 5500 10532
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 6368 10412 6420 10464
rect 8116 10616 8168 10668
rect 7932 10548 7984 10600
rect 9496 10684 9548 10736
rect 9128 10616 9180 10668
rect 9312 10616 9364 10668
rect 11520 10727 11572 10736
rect 11520 10693 11529 10727
rect 11529 10693 11563 10727
rect 11563 10693 11572 10727
rect 11520 10684 11572 10693
rect 17040 10752 17092 10804
rect 12440 10727 12492 10736
rect 12440 10693 12449 10727
rect 12449 10693 12483 10727
rect 12483 10693 12492 10727
rect 12440 10684 12492 10693
rect 15476 10684 15528 10736
rect 15936 10684 15988 10736
rect 16212 10684 16264 10736
rect 16948 10727 17000 10736
rect 16948 10693 16957 10727
rect 16957 10693 16991 10727
rect 16991 10693 17000 10727
rect 16948 10684 17000 10693
rect 8576 10480 8628 10532
rect 8668 10412 8720 10464
rect 11060 10480 11112 10532
rect 13268 10616 13320 10668
rect 15660 10616 15712 10668
rect 12256 10548 12308 10600
rect 14740 10548 14792 10600
rect 13084 10412 13136 10464
rect 14464 10412 14516 10464
rect 17868 10412 17920 10464
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 4436 10208 4488 10260
rect 14924 10208 14976 10260
rect 15844 10208 15896 10260
rect 2320 10140 2372 10192
rect 6000 10140 6052 10192
rect 3240 9868 3292 9920
rect 3700 9868 3752 9920
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 11796 10140 11848 10192
rect 16212 10140 16264 10192
rect 8024 10072 8076 10124
rect 9128 10072 9180 10124
rect 10324 10072 10376 10124
rect 10876 10072 10928 10124
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 12348 10072 12400 10124
rect 17960 10072 18012 10124
rect 18420 10072 18472 10124
rect 10600 10004 10652 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 8208 9936 8260 9988
rect 8576 9936 8628 9988
rect 8668 9979 8720 9988
rect 8668 9945 8677 9979
rect 8677 9945 8711 9979
rect 8711 9945 8720 9979
rect 8668 9936 8720 9945
rect 11520 9936 11572 9988
rect 10324 9868 10376 9920
rect 10692 9868 10744 9920
rect 10784 9868 10836 9920
rect 12256 9868 12308 9920
rect 15936 9868 15988 9920
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 7012 9664 7064 9716
rect 8484 9664 8536 9716
rect 12624 9664 12676 9716
rect 12992 9664 13044 9716
rect 16856 9664 16908 9716
rect 4252 9596 4304 9648
rect 5540 9596 5592 9648
rect 8944 9596 8996 9648
rect 9404 9639 9456 9648
rect 9404 9605 9413 9639
rect 9413 9605 9447 9639
rect 9447 9605 9456 9639
rect 9404 9596 9456 9605
rect 9772 9596 9824 9648
rect 10784 9596 10836 9648
rect 13820 9596 13872 9648
rect 14556 9596 14608 9648
rect 6368 9528 6420 9580
rect 1676 9460 1728 9512
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7288 9528 7340 9580
rect 7748 9528 7800 9580
rect 10048 9571 10100 9580
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 7564 9460 7616 9512
rect 5540 9392 5592 9444
rect 6736 9392 6788 9444
rect 9404 9460 9456 9512
rect 5908 9324 5960 9376
rect 7012 9324 7064 9376
rect 8208 9392 8260 9444
rect 11796 9460 11848 9512
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 13084 9528 13136 9580
rect 13176 9528 13228 9580
rect 15476 9528 15528 9580
rect 15844 9528 15896 9580
rect 16396 9528 16448 9580
rect 7840 9324 7892 9376
rect 8392 9324 8444 9376
rect 10968 9324 11020 9376
rect 16856 9392 16908 9444
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 3792 9120 3844 9172
rect 6092 9120 6144 9172
rect 5356 9052 5408 9104
rect 7288 9120 7340 9172
rect 7564 9052 7616 9104
rect 7840 9052 7892 9104
rect 8116 9052 8168 9104
rect 4712 8984 4764 9036
rect 9128 9052 9180 9104
rect 10416 9120 10468 9172
rect 10508 9120 10560 9172
rect 11060 9120 11112 9172
rect 11980 9120 12032 9172
rect 13912 9120 13964 9172
rect 4436 8916 4488 8968
rect 6092 8916 6144 8968
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7656 8916 7708 8968
rect 8024 8916 8076 8968
rect 8668 8916 8720 8968
rect 9496 8984 9548 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9772 8984 9824 9036
rect 10140 8984 10192 9036
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 10692 9052 10744 9104
rect 11796 8984 11848 9036
rect 13452 9052 13504 9104
rect 15568 9052 15620 9104
rect 15936 9052 15988 9104
rect 15292 8984 15344 9036
rect 2412 8848 2464 8900
rect 4988 8848 5040 8900
rect 5540 8848 5592 8900
rect 6736 8848 6788 8900
rect 4068 8780 4120 8832
rect 6368 8780 6420 8832
rect 7288 8848 7340 8900
rect 9404 8848 9456 8900
rect 7104 8780 7156 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 9312 8780 9364 8832
rect 10048 8780 10100 8832
rect 10692 8891 10744 8900
rect 10692 8857 10701 8891
rect 10701 8857 10735 8891
rect 10735 8857 10744 8891
rect 10692 8848 10744 8857
rect 13912 8916 13964 8968
rect 14280 8916 14332 8968
rect 11428 8848 11480 8900
rect 11888 8848 11940 8900
rect 12256 8891 12308 8900
rect 12256 8857 12265 8891
rect 12265 8857 12299 8891
rect 12299 8857 12308 8891
rect 12256 8848 12308 8857
rect 18696 8848 18748 8900
rect 11152 8780 11204 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 3792 8576 3844 8628
rect 4160 8576 4212 8628
rect 5172 8576 5224 8628
rect 6000 8576 6052 8628
rect 9496 8576 9548 8628
rect 9588 8576 9640 8628
rect 10784 8576 10836 8628
rect 11428 8576 11480 8628
rect 12992 8576 13044 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 14096 8576 14148 8628
rect 14188 8619 14240 8628
rect 14188 8585 14197 8619
rect 14197 8585 14231 8619
rect 14231 8585 14240 8619
rect 14188 8576 14240 8585
rect 14372 8576 14424 8628
rect 3516 8508 3568 8560
rect 5448 8508 5500 8560
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 3516 8372 3568 8424
rect 4160 8440 4212 8492
rect 5632 8440 5684 8492
rect 6092 8440 6144 8492
rect 6276 8508 6328 8560
rect 6368 8372 6420 8424
rect 6828 8440 6880 8492
rect 7656 8440 7708 8492
rect 8116 8508 8168 8560
rect 9404 8440 9456 8492
rect 10416 8508 10468 8560
rect 10876 8508 10928 8560
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 12164 8508 12216 8517
rect 12348 8551 12400 8560
rect 12348 8517 12357 8551
rect 12357 8517 12391 8551
rect 12391 8517 12400 8551
rect 12348 8508 12400 8517
rect 6920 8372 6972 8424
rect 7104 8372 7156 8424
rect 7748 8372 7800 8424
rect 8024 8372 8076 8424
rect 9680 8372 9732 8424
rect 7840 8304 7892 8356
rect 7932 8304 7984 8356
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 9220 8304 9272 8356
rect 9496 8304 9548 8356
rect 4528 8236 4580 8288
rect 9680 8236 9732 8288
rect 9956 8304 10008 8356
rect 10140 8254 10192 8306
rect 10232 8347 10284 8356
rect 10232 8313 10241 8347
rect 10241 8313 10275 8347
rect 10275 8313 10284 8347
rect 10232 8304 10284 8313
rect 10416 8304 10468 8356
rect 10876 8347 10928 8356
rect 10876 8313 10885 8347
rect 10885 8313 10919 8347
rect 10919 8313 10928 8347
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13820 8440 13872 8492
rect 11888 8372 11940 8424
rect 10876 8304 10928 8313
rect 13084 8372 13136 8424
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14740 8440 14792 8492
rect 13176 8304 13228 8356
rect 13452 8304 13504 8356
rect 18512 8236 18564 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 3332 8032 3384 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 6184 7964 6236 8016
rect 11060 7964 11112 8016
rect 1768 7760 1820 7812
rect 2320 7760 2372 7812
rect 2964 7828 3016 7880
rect 4436 7896 4488 7948
rect 8116 7896 8168 7948
rect 8760 7896 8812 7948
rect 9588 7896 9640 7948
rect 9956 7896 10008 7948
rect 3424 7760 3476 7812
rect 4252 7828 4304 7880
rect 4160 7692 4212 7744
rect 5080 7803 5132 7812
rect 5080 7769 5089 7803
rect 5089 7769 5123 7803
rect 5123 7769 5132 7803
rect 5080 7760 5132 7769
rect 5540 7760 5592 7812
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 7656 7828 7708 7880
rect 8300 7828 8352 7880
rect 10140 7828 10192 7880
rect 10416 7828 10468 7880
rect 10508 7828 10560 7880
rect 10876 7828 10928 7880
rect 11612 8032 11664 8084
rect 12900 8032 12952 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 13728 8032 13780 8084
rect 13820 8032 13872 8084
rect 15016 8032 15068 8084
rect 11796 7896 11848 7948
rect 15292 7964 15344 8016
rect 5724 7692 5776 7744
rect 6368 7692 6420 7744
rect 6920 7692 6972 7744
rect 7748 7692 7800 7744
rect 8116 7692 8168 7744
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 12716 7760 12768 7812
rect 11888 7692 11940 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 13728 7896 13780 7948
rect 13912 7828 13964 7880
rect 15016 7828 15068 7880
rect 15752 7828 15804 7880
rect 18144 7828 18196 7880
rect 16672 7760 16724 7812
rect 16948 7760 17000 7812
rect 12900 7692 12952 7701
rect 14188 7692 14240 7744
rect 14648 7692 14700 7744
rect 16580 7692 16632 7744
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 1768 7488 1820 7540
rect 2228 7488 2280 7540
rect 2596 7420 2648 7472
rect 3148 7420 3200 7472
rect 6828 7488 6880 7540
rect 7472 7488 7524 7540
rect 10324 7531 10376 7540
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 1676 7284 1728 7336
rect 3424 7284 3476 7336
rect 6276 7420 6328 7472
rect 10508 7420 10560 7472
rect 4252 7284 4304 7336
rect 5356 7284 5408 7336
rect 5724 7284 5776 7336
rect 7104 7352 7156 7404
rect 7840 7352 7892 7404
rect 10324 7352 10376 7404
rect 10692 7352 10744 7404
rect 11796 7488 11848 7540
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 15292 7488 15344 7540
rect 10968 7463 11020 7472
rect 10968 7429 10977 7463
rect 10977 7429 11011 7463
rect 11011 7429 11020 7463
rect 10968 7420 11020 7429
rect 11520 7463 11572 7472
rect 11520 7429 11529 7463
rect 11529 7429 11563 7463
rect 11563 7429 11572 7463
rect 11520 7420 11572 7429
rect 13636 7420 13688 7472
rect 15108 7420 15160 7472
rect 15384 7420 15436 7472
rect 13360 7352 13412 7404
rect 17316 7488 17368 7540
rect 6092 7284 6144 7336
rect 2320 7148 2372 7200
rect 2504 7148 2556 7200
rect 3700 7148 3752 7200
rect 10784 7284 10836 7336
rect 14004 7284 14056 7336
rect 15108 7284 15160 7336
rect 16948 7352 17000 7404
rect 7104 7216 7156 7268
rect 12808 7216 12860 7268
rect 13820 7216 13872 7268
rect 14372 7216 14424 7268
rect 14832 7216 14884 7268
rect 15660 7216 15712 7268
rect 15936 7216 15988 7268
rect 16120 7216 16172 7268
rect 7012 7148 7064 7200
rect 7472 7148 7524 7200
rect 7840 7148 7892 7200
rect 11336 7148 11388 7200
rect 12348 7148 12400 7200
rect 13452 7148 13504 7200
rect 13636 7148 13688 7200
rect 16304 7148 16356 7200
rect 17960 7259 18012 7268
rect 17960 7225 17969 7259
rect 17969 7225 18003 7259
rect 18003 7225 18012 7259
rect 17960 7216 18012 7225
rect 17592 7191 17644 7200
rect 17592 7157 17601 7191
rect 17601 7157 17635 7191
rect 17635 7157 17644 7191
rect 17592 7148 17644 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 2320 6944 2372 6996
rect 2688 6944 2740 6996
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5816 6944 5868 6996
rect 7840 6944 7892 6996
rect 8576 6944 8628 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 9588 6944 9640 6996
rect 6368 6876 6420 6928
rect 3516 6808 3568 6860
rect 4252 6808 4304 6860
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 10600 6876 10652 6928
rect 10692 6876 10744 6928
rect 10968 6876 11020 6928
rect 12164 6944 12216 6996
rect 12532 6944 12584 6996
rect 12624 6987 12676 6996
rect 12624 6953 12633 6987
rect 12633 6953 12667 6987
rect 12667 6953 12676 6987
rect 12624 6944 12676 6953
rect 14004 6944 14056 6996
rect 17592 6944 17644 6996
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 18144 6944 18196 6996
rect 9312 6808 9364 6860
rect 3976 6672 4028 6724
rect 4804 6672 4856 6724
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 9128 6740 9180 6792
rect 9496 6808 9548 6860
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 14648 6876 14700 6928
rect 14924 6876 14976 6928
rect 15384 6876 15436 6928
rect 11336 6783 11388 6792
rect 11336 6749 11337 6783
rect 11337 6749 11371 6783
rect 11371 6749 11388 6783
rect 11336 6740 11388 6749
rect 8944 6672 8996 6724
rect 9496 6715 9548 6724
rect 9496 6681 9505 6715
rect 9505 6681 9539 6715
rect 9539 6681 9548 6715
rect 9496 6672 9548 6681
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 12348 6808 12400 6860
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 12440 6740 12492 6792
rect 13912 6808 13964 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 14740 6808 14792 6860
rect 14832 6740 14884 6792
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15108 6740 15160 6792
rect 15752 6740 15804 6792
rect 16028 6740 16080 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 2504 6604 2556 6656
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3792 6604 3844 6656
rect 5724 6604 5776 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 7472 6604 7524 6656
rect 8576 6604 8628 6656
rect 10600 6604 10652 6656
rect 11336 6604 11388 6656
rect 12256 6715 12308 6724
rect 12256 6681 12265 6715
rect 12265 6681 12299 6715
rect 12299 6681 12308 6715
rect 12256 6672 12308 6681
rect 11704 6604 11756 6656
rect 11980 6604 12032 6656
rect 12164 6604 12216 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 13820 6672 13872 6724
rect 14372 6672 14424 6724
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 13636 6604 13688 6656
rect 14648 6604 14700 6656
rect 17132 6672 17184 6724
rect 16028 6604 16080 6656
rect 18512 6672 18564 6724
rect 18052 6604 18104 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 5632 6400 5684 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 10232 6400 10284 6452
rect 11888 6443 11940 6452
rect 11888 6409 11913 6443
rect 11913 6409 11940 6443
rect 11888 6400 11940 6409
rect 12164 6400 12216 6452
rect 13912 6400 13964 6452
rect 14096 6400 14148 6452
rect 15200 6400 15252 6452
rect 17316 6443 17368 6452
rect 17316 6409 17325 6443
rect 17325 6409 17359 6443
rect 17359 6409 17368 6443
rect 17316 6400 17368 6409
rect 3056 6332 3108 6384
rect 3792 6264 3844 6316
rect 4436 6264 4488 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 6644 6264 6696 6316
rect 7012 6332 7064 6384
rect 9680 6332 9732 6384
rect 11704 6375 11756 6384
rect 11704 6341 11713 6375
rect 11713 6341 11747 6375
rect 11747 6341 11756 6375
rect 11704 6332 11756 6341
rect 10784 6264 10836 6316
rect 11060 6264 11112 6316
rect 14280 6332 14332 6384
rect 15108 6332 15160 6384
rect 16120 6332 16172 6384
rect 16580 6332 16632 6384
rect 12900 6264 12952 6316
rect 15292 6264 15344 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 16672 6264 16724 6316
rect 17132 6375 17184 6384
rect 17132 6341 17141 6375
rect 17141 6341 17175 6375
rect 17175 6341 17184 6375
rect 17132 6332 17184 6341
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17408 6332 17460 6384
rect 17500 6264 17552 6316
rect 18144 6307 18196 6316
rect 18144 6273 18153 6307
rect 18153 6273 18187 6307
rect 18187 6273 18196 6307
rect 18144 6264 18196 6273
rect 18236 6264 18288 6316
rect 4804 6196 4856 6248
rect 8852 6196 8904 6248
rect 8944 6196 8996 6248
rect 10508 6196 10560 6248
rect 10600 6196 10652 6248
rect 11704 6196 11756 6248
rect 4252 6128 4304 6180
rect 7472 6128 7524 6180
rect 4528 6060 4580 6112
rect 6000 6060 6052 6112
rect 6828 6060 6880 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 13820 6196 13872 6248
rect 12164 6128 12216 6180
rect 12624 6128 12676 6180
rect 12716 6128 12768 6180
rect 13084 6128 13136 6180
rect 16672 6128 16724 6180
rect 16856 6171 16908 6180
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 17776 6196 17828 6248
rect 11336 6060 11388 6069
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 12256 6060 12308 6112
rect 12532 6060 12584 6112
rect 13820 6060 13872 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 3240 5856 3292 5908
rect 3700 5856 3752 5908
rect 4620 5856 4672 5908
rect 4436 5788 4488 5840
rect 7380 5856 7432 5908
rect 9772 5856 9824 5908
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 12532 5856 12584 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 4804 5788 4856 5840
rect 5448 5788 5500 5840
rect 5724 5788 5776 5840
rect 3148 5763 3200 5772
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 4068 5652 4120 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 10876 5788 10928 5840
rect 15108 5856 15160 5908
rect 15292 5856 15344 5908
rect 13360 5788 13412 5840
rect 13636 5788 13688 5840
rect 17224 5856 17276 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 18236 5856 18288 5908
rect 9496 5720 9548 5772
rect 12624 5720 12676 5772
rect 9772 5652 9824 5704
rect 10048 5652 10100 5704
rect 14372 5720 14424 5772
rect 15660 5720 15712 5772
rect 16580 5720 16632 5772
rect 12900 5652 12952 5704
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 17500 5652 17552 5704
rect 6368 5584 6420 5636
rect 8300 5584 8352 5636
rect 9588 5584 9640 5636
rect 10600 5627 10652 5636
rect 10600 5593 10609 5627
rect 10609 5593 10643 5627
rect 10643 5593 10652 5627
rect 10600 5584 10652 5593
rect 10784 5627 10836 5636
rect 10784 5593 10809 5627
rect 10809 5593 10836 5627
rect 10784 5584 10836 5593
rect 4068 5516 4120 5568
rect 4252 5516 4304 5568
rect 4436 5559 4488 5568
rect 4436 5525 4445 5559
rect 4445 5525 4479 5559
rect 4479 5525 4488 5559
rect 4436 5516 4488 5525
rect 10508 5516 10560 5568
rect 12808 5584 12860 5636
rect 13084 5584 13136 5636
rect 13268 5627 13320 5636
rect 13268 5593 13295 5627
rect 13295 5593 13320 5627
rect 13268 5584 13320 5593
rect 13360 5584 13412 5636
rect 13820 5584 13872 5636
rect 15752 5584 15804 5636
rect 17132 5584 17184 5636
rect 17776 5584 17828 5636
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 1584 5312 1636 5364
rect 7380 5312 7432 5364
rect 2412 5287 2464 5296
rect 2412 5253 2421 5287
rect 2421 5253 2455 5287
rect 2455 5253 2464 5287
rect 2412 5244 2464 5253
rect 4436 5244 4488 5296
rect 9312 5312 9364 5364
rect 9588 5312 9640 5364
rect 10784 5312 10836 5364
rect 13084 5312 13136 5364
rect 13820 5312 13872 5364
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 2504 5176 2556 5228
rect 5816 5176 5868 5228
rect 8208 5244 8260 5296
rect 9036 5244 9088 5296
rect 9956 5244 10008 5296
rect 11612 5244 11664 5296
rect 7564 5176 7616 5228
rect 1860 5108 1912 5160
rect 4252 5108 4304 5160
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 10324 5176 10376 5228
rect 15936 5176 15988 5228
rect 11336 5108 11388 5160
rect 16764 5312 16816 5364
rect 16488 5244 16540 5296
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 18052 5312 18104 5364
rect 16580 5176 16632 5228
rect 17500 5176 17552 5228
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 17132 5108 17184 5160
rect 9312 5040 9364 5092
rect 6828 4972 6880 5024
rect 9956 4972 10008 5024
rect 10140 5083 10192 5092
rect 10140 5049 10149 5083
rect 10149 5049 10183 5083
rect 10183 5049 10192 5083
rect 10140 5040 10192 5049
rect 10324 5040 10376 5092
rect 16580 5040 16632 5092
rect 13084 4972 13136 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 15476 4972 15528 5024
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 16948 4972 17000 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 1768 4768 1820 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 4988 4768 5040 4820
rect 6828 4768 6880 4820
rect 7288 4768 7340 4820
rect 7564 4768 7616 4820
rect 8484 4768 8536 4820
rect 10324 4768 10376 4820
rect 10600 4768 10652 4820
rect 13084 4768 13136 4820
rect 15200 4768 15252 4820
rect 16488 4768 16540 4820
rect 16580 4811 16632 4820
rect 16580 4777 16589 4811
rect 16589 4777 16623 4811
rect 16623 4777 16632 4811
rect 16580 4768 16632 4777
rect 16856 4768 16908 4820
rect 7380 4700 7432 4752
rect 8576 4700 8628 4752
rect 10416 4700 10468 4752
rect 10692 4700 10744 4752
rect 11152 4700 11204 4752
rect 6092 4632 6144 4684
rect 8300 4632 8352 4684
rect 4344 4564 4396 4616
rect 6184 4564 6236 4616
rect 6828 4564 6880 4616
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 5816 4496 5868 4548
rect 9588 4564 9640 4616
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 11152 4539 11204 4548
rect 11152 4505 11161 4539
rect 11161 4505 11195 4539
rect 11195 4505 11204 4539
rect 11152 4496 11204 4505
rect 10876 4428 10928 4480
rect 15108 4700 15160 4752
rect 15292 4700 15344 4752
rect 13452 4632 13504 4684
rect 13268 4564 13320 4616
rect 18328 4768 18380 4820
rect 18696 4700 18748 4752
rect 14924 4539 14976 4548
rect 14924 4505 14933 4539
rect 14933 4505 14967 4539
rect 14967 4505 14976 4539
rect 14924 4496 14976 4505
rect 15108 4539 15160 4548
rect 15108 4505 15117 4539
rect 15117 4505 15151 4539
rect 15151 4505 15160 4539
rect 15108 4496 15160 4505
rect 15292 4539 15344 4548
rect 15292 4505 15301 4539
rect 15301 4505 15335 4539
rect 15335 4505 15344 4539
rect 15292 4496 15344 4505
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 18144 4496 18196 4548
rect 15016 4428 15068 4480
rect 18420 4471 18472 4480
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 3884 4224 3936 4276
rect 4068 4224 4120 4276
rect 6368 4224 6420 4276
rect 7380 4267 7432 4276
rect 7380 4233 7389 4267
rect 7389 4233 7423 4267
rect 7423 4233 7432 4267
rect 7380 4224 7432 4233
rect 8484 4224 8536 4276
rect 8668 4267 8720 4276
rect 8668 4233 8695 4267
rect 8695 4233 8720 4267
rect 8668 4224 8720 4233
rect 11060 4224 11112 4276
rect 2504 4156 2556 4208
rect 4252 4199 4304 4208
rect 4252 4165 4261 4199
rect 4261 4165 4295 4199
rect 4295 4165 4304 4199
rect 4252 4156 4304 4165
rect 8300 4156 8352 4208
rect 8944 4156 8996 4208
rect 9036 4156 9088 4208
rect 9680 4156 9732 4208
rect 10048 4156 10100 4208
rect 11152 4156 11204 4208
rect 11612 4156 11664 4208
rect 14004 4224 14056 4276
rect 15568 4224 15620 4276
rect 13728 4156 13780 4208
rect 18144 4156 18196 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6736 4088 6788 4140
rect 3516 4020 3568 4072
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 4620 4020 4672 4072
rect 8208 3952 8260 4004
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 6828 3884 6880 3936
rect 8116 3884 8168 3936
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 11244 4020 11296 4072
rect 11796 4020 11848 4072
rect 18696 4088 18748 4140
rect 14832 4020 14884 4072
rect 16672 3952 16724 4004
rect 9588 3884 9640 3936
rect 10232 3884 10284 3936
rect 13544 3884 13596 3936
rect 17868 3927 17920 3936
rect 17868 3893 17877 3927
rect 17877 3893 17911 3927
rect 17911 3893 17920 3927
rect 17868 3884 17920 3893
rect 18144 3884 18196 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 1860 3680 1912 3732
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 5540 3680 5592 3732
rect 6460 3680 6512 3732
rect 12072 3680 12124 3732
rect 16396 3680 16448 3732
rect 9496 3612 9548 3664
rect 11336 3655 11388 3664
rect 11336 3621 11345 3655
rect 11345 3621 11379 3655
rect 11379 3621 11388 3655
rect 11336 3612 11388 3621
rect 13820 3612 13872 3664
rect 3976 3544 4028 3596
rect 8024 3544 8076 3596
rect 9220 3544 9272 3596
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 9956 3544 10008 3596
rect 2964 3476 3016 3528
rect 9496 3476 9548 3528
rect 10968 3476 11020 3528
rect 5264 3408 5316 3460
rect 8668 3408 8720 3460
rect 8944 3451 8996 3460
rect 8944 3417 8953 3451
rect 8953 3417 8987 3451
rect 8987 3417 8996 3451
rect 8944 3408 8996 3417
rect 9036 3408 9088 3460
rect 4160 3340 4212 3392
rect 9956 3408 10008 3460
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3340 9456 3392
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 18788 3476 18840 3528
rect 11520 3340 11572 3392
rect 17316 3408 17368 3460
rect 12164 3340 12216 3392
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 16212 3340 16264 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 1768 3136 1820 3188
rect 10048 3136 10100 3188
rect 10876 3136 10928 3188
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 14372 3136 14424 3188
rect 15108 3136 15160 3188
rect 15752 3136 15804 3188
rect 8944 3068 8996 3120
rect 10508 3068 10560 3120
rect 11520 3111 11572 3120
rect 11520 3077 11529 3111
rect 11529 3077 11563 3111
rect 11563 3077 11572 3111
rect 11520 3068 11572 3077
rect 8668 3000 8720 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12072 3068 12124 3120
rect 12440 3068 12492 3120
rect 12992 3000 13044 3052
rect 5540 2796 5592 2848
rect 11888 2864 11940 2916
rect 12164 2864 12216 2916
rect 17408 2864 17460 2916
rect 6828 2796 6880 2848
rect 8392 2796 8444 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 11428 2592 11480 2644
rect 15200 2592 15252 2644
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 11704 2524 11756 2576
rect 14924 2567 14976 2576
rect 14924 2533 14933 2567
rect 14933 2533 14967 2567
rect 14967 2533 14976 2567
rect 14924 2524 14976 2533
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 16120 2456 16172 2508
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 3608 2320 3660 2372
rect 13176 2320 13228 2372
rect 14372 2320 14424 2372
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 18604 2388 18656 2440
rect 11796 2252 11848 2304
rect 18420 2295 18472 2304
rect 18420 2261 18429 2295
rect 18429 2261 18463 2295
rect 18463 2261 18472 2295
rect 18420 2252 18472 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
<< metal2 >>
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 7300 17134 7328 17546
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1676 16584 1728 16590
rect 1780 16574 1808 16730
rect 3160 16726 3188 16934
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3330 16688 3386 16697
rect 1780 16546 1900 16574
rect 1676 16526 1728 16532
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15094 1624 15438
rect 1584 15088 1636 15094
rect 1582 15056 1584 15065
rect 1636 15056 1638 15065
rect 1582 14991 1638 15000
rect 1688 14414 1716 16526
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1398 13424 1454 13433
rect 1398 13359 1454 13368
rect 1412 4049 1440 13359
rect 1582 12744 1638 12753
rect 1582 12679 1638 12688
rect 1596 5370 1624 12679
rect 1688 9625 1716 14350
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 8430 1716 9454
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7342 1716 8366
rect 1780 7818 1808 12718
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1780 4826 1808 7482
rect 1872 5166 1900 16546
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15337 2176 15370
rect 2412 15360 2464 15366
rect 2134 15328 2190 15337
rect 2412 15302 2464 15308
rect 2134 15263 2190 15272
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 2332 14414 2360 14758
rect 2424 14414 2452 15302
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2240 11762 2268 12378
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 2332 10810 2360 14214
rect 2424 13870 2452 14350
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11898 2452 12038
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1952 8424 2004 8430
rect 1950 8392 1952 8401
rect 2004 8392 2006 8401
rect 1950 8327 2006 8336
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2332 7970 2360 10134
rect 2424 9489 2452 11698
rect 2516 10674 2544 15506
rect 3160 15348 3188 16662
rect 3330 16623 3386 16632
rect 3160 15320 3280 15348
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 3146 15192 3202 15201
rect 3146 15127 3202 15136
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 13297 2636 13806
rect 2594 13288 2650 13297
rect 2594 13223 2650 13232
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2594 10704 2650 10713
rect 2504 10668 2556 10674
rect 2594 10639 2650 10648
rect 2504 10610 2556 10616
rect 2608 10554 2636 10639
rect 2516 10526 2636 10554
rect 2410 9480 2466 9489
rect 2410 9415 2466 9424
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2240 7942 2360 7970
rect 2240 7546 2268 7942
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2332 7206 2360 7754
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5710 2360 6938
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2424 5302 2452 8842
rect 2516 7426 2544 10526
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2976 7886 3004 12786
rect 3054 12744 3110 12753
rect 3054 12679 3056 12688
rect 3108 12679 3110 12688
rect 3056 12650 3108 12656
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3068 11558 3096 11698
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3054 9752 3110 9761
rect 3054 9687 3110 9696
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2596 7472 2648 7478
rect 2516 7420 2596 7426
rect 2516 7414 2648 7420
rect 2686 7440 2742 7449
rect 2516 7398 2636 7414
rect 2686 7375 2742 7384
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2516 6662 2544 7142
rect 2700 7002 2728 7375
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 2516 4214 2544 5170
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3194 1808 3878
rect 1872 3738 1900 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2976 3738 3004 7822
rect 3068 7449 3096 9687
rect 3160 7478 3188 15127
rect 3252 9926 3280 15320
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 7472 3200 7478
rect 3054 7440 3110 7449
rect 3148 7414 3200 7420
rect 3054 7375 3110 7384
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6390 3096 6598
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3160 5778 3188 6287
rect 3252 5914 3280 9454
rect 3344 8090 3372 16623
rect 3436 8090 3464 17002
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16794 4292 16934
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3804 16590 3832 16662
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3804 15910 3832 16526
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3528 13938 3556 14554
rect 3804 14414 3832 15846
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 12442 3556 12786
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3528 8566 3556 12242
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 8265 3556 8366
rect 3514 8256 3570 8265
rect 3514 8191 3570 8200
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3424 7812 3476 7818
rect 3476 7772 3556 7800
rect 3424 7754 3476 7760
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 6848 3464 7278
rect 3528 7041 3556 7772
rect 3514 7032 3570 7041
rect 3514 6967 3516 6976
rect 3568 6967 3570 6976
rect 3516 6938 3568 6944
rect 3516 6860 3568 6866
rect 3436 6820 3516 6848
rect 3516 6802 3568 6808
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3528 4078 3556 6802
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2976 3534 3004 3674
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3620 2378 3648 13126
rect 3698 13016 3754 13025
rect 3698 12951 3754 12960
rect 3712 12918 3740 12951
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3804 12850 3832 14350
rect 3896 13326 3924 15574
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 14006 4108 15302
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4068 14000 4120 14006
rect 4066 13968 4068 13977
rect 4120 13968 4122 13977
rect 4066 13903 4122 13912
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3804 11830 3832 12106
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3700 11552 3752 11558
rect 3698 11520 3700 11529
rect 3752 11520 3754 11529
rect 3698 11455 3754 11464
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 7206 3740 9862
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3804 8634 3832 9114
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3896 7993 3924 12174
rect 3976 12096 4028 12102
rect 4080 12084 4108 12650
rect 4028 12056 4108 12084
rect 3976 12038 4028 12044
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3882 7984 3938 7993
rect 3882 7919 3938 7928
rect 3882 7848 3938 7857
rect 3882 7783 3938 7792
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 5914 3740 7142
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6458 3832 6598
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3804 6322 3832 6394
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3896 4282 3924 7783
rect 3988 6730 4016 11562
rect 4080 10577 4108 12056
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4080 9092 4108 10503
rect 4172 9194 4200 14826
rect 4264 9654 4292 16390
rect 4356 14618 4384 16458
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4894 15464 4950 15473
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4356 12238 4384 14554
rect 4448 13530 4476 15438
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4434 13424 4490 13433
rect 4434 13359 4490 13368
rect 4448 13326 4476 13359
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4356 12102 4384 12174
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 10169 4384 12038
rect 4448 11218 4476 12310
rect 4526 11792 4582 11801
rect 4526 11727 4528 11736
rect 4580 11727 4582 11736
rect 4528 11698 4580 11704
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 10266 4476 10406
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4526 9616 4582 9625
rect 4526 9551 4582 9560
rect 4172 9166 4292 9194
rect 4080 9064 4200 9092
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4080 8838 4108 8871
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4066 8664 4122 8673
rect 4172 8634 4200 9064
rect 4264 8673 4292 9166
rect 4342 9072 4398 9081
rect 4342 9007 4398 9016
rect 4250 8664 4306 8673
rect 4066 8599 4122 8608
rect 4160 8628 4212 8634
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4080 5710 4108 8599
rect 4250 8599 4306 8608
rect 4160 8570 4212 8576
rect 4158 8528 4214 8537
rect 4158 8463 4160 8472
rect 4212 8463 4214 8472
rect 4160 8434 4212 8440
rect 4250 8392 4306 8401
rect 4250 8327 4306 8336
rect 4264 8022 4292 8327
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 4282 4108 5510
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3602 4016 4014
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4172 3398 4200 7686
rect 4264 7342 4292 7822
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4264 6866 4292 7278
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4264 5574 4292 6122
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4264 4214 4292 5102
rect 4356 4826 4384 9007
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4448 7954 4476 8910
rect 4540 8294 4568 9551
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4540 6322 4568 8230
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4448 5846 4476 6258
rect 4540 6118 4568 6258
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4632 5914 4660 15438
rect 4712 15428 4764 15434
rect 4894 15399 4896 15408
rect 4712 15370 4764 15376
rect 4948 15399 4950 15408
rect 4896 15370 4948 15376
rect 4724 12209 4752 15370
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 14074 4936 14350
rect 5000 14074 5028 16390
rect 5092 14482 5120 16594
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 15366 5304 16526
rect 6092 16516 6144 16522
rect 6092 16458 6144 16464
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 5460 15502 5488 15535
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5092 13870 5120 14282
rect 5184 14006 5212 14418
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 13394 4936 13670
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4710 12200 4766 12209
rect 4710 12135 4766 12144
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11830 4844 12038
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4816 10810 4844 11766
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5302 4476 5510
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4356 4622 4384 4762
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4632 4078 4660 5850
rect 4724 5710 4752 8978
rect 4816 8401 4844 10746
rect 4802 8392 4858 8401
rect 4802 8327 4858 8336
rect 4802 6760 4858 6769
rect 4802 6695 4804 6704
rect 4856 6695 4858 6704
rect 4804 6666 4856 6672
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5846 4844 6190
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4804 5704 4856 5710
rect 4908 5692 4936 13330
rect 5000 11626 5028 13466
rect 5092 12434 5120 13806
rect 5184 13258 5212 13806
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5276 12434 5304 15302
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5092 12406 5212 12434
rect 5276 12406 5396 12434
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4856 5664 4936 5692
rect 4804 5646 4856 5652
rect 5000 4826 5028 8842
rect 5092 7818 5120 11222
rect 5184 8634 5212 12406
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 5276 3466 5304 11222
rect 5368 9110 5396 12406
rect 5460 12102 5488 13466
rect 5552 13138 5580 13942
rect 5644 13569 5672 16390
rect 5828 16238 6040 16266
rect 5828 16182 5856 16238
rect 6012 16182 6040 16238
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5724 15496 5776 15502
rect 5828 15484 5856 15846
rect 5776 15456 5856 15484
rect 5724 15438 5776 15444
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5736 14890 5764 14962
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5630 13560 5686 13569
rect 5630 13495 5686 13504
rect 5552 13110 5672 13138
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8401 5396 9046
rect 5460 8566 5488 10474
rect 5552 9654 5580 12582
rect 5644 11665 5672 13110
rect 5630 11656 5686 11665
rect 5630 11591 5686 11600
rect 5736 10010 5764 14486
rect 5644 9982 5764 10010
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 8906 5580 9386
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5644 8498 5672 9982
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5354 8392 5410 8401
rect 5354 8327 5410 8336
rect 5736 8265 5764 9862
rect 5722 8256 5778 8265
rect 5722 8191 5778 8200
rect 5828 7936 5856 15456
rect 5920 10742 5948 16118
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 6012 14550 6040 15370
rect 6104 15337 6132 16458
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15570 6224 15982
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6090 15328 6146 15337
rect 6090 15263 6146 15272
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 14006 6040 14214
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 12714 6040 13670
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 6012 10198 6040 12378
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5998 9616 6054 9625
rect 5998 9551 6054 9560
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5460 7908 5856 7936
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5368 6225 5396 7278
rect 5354 6216 5410 6225
rect 5354 6151 5410 6160
rect 5354 6080 5410 6089
rect 5354 6015 5410 6024
rect 5368 3641 5396 6015
rect 5460 5846 5488 7908
rect 5920 7857 5948 9318
rect 6012 8809 6040 9551
rect 6104 9178 6132 15030
rect 6196 14822 6224 15506
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 13938 6224 14758
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6196 13394 6224 13874
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12918 6224 13330
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6196 12306 6224 12854
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11762 6224 12242
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6104 8974 6132 9114
rect 6092 8968 6144 8974
rect 6288 8945 6316 16390
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6380 15706 6408 15982
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6366 15600 6422 15609
rect 7300 15570 7328 17070
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 6366 15535 6368 15544
rect 6420 15535 6422 15544
rect 6644 15564 6696 15570
rect 6368 15506 6420 15512
rect 6644 15506 6696 15512
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6380 12646 6408 14826
rect 6472 14618 6500 15030
rect 6656 14618 6684 15506
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 7300 14074 7328 15506
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6472 13734 6500 13942
rect 6748 13841 6776 14010
rect 6734 13832 6790 13841
rect 6734 13767 6790 13776
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6472 12186 6500 13194
rect 6564 13161 6592 13670
rect 6656 13190 6684 13670
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6644 13184 6696 13190
rect 6550 13152 6606 13161
rect 6644 13126 6696 13132
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6550 13087 6606 13096
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6472 12158 6592 12186
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 9761 6408 10406
rect 6366 9752 6422 9761
rect 6366 9687 6422 9696
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6092 8910 6144 8916
rect 6274 8936 6330 8945
rect 6274 8871 6330 8880
rect 6380 8838 6408 9522
rect 6368 8832 6420 8838
rect 5998 8800 6054 8809
rect 5998 8735 6054 8744
rect 6274 8800 6330 8809
rect 6368 8774 6420 8780
rect 6274 8735 6330 8744
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5906 7848 5962 7857
rect 5540 7812 5592 7818
rect 5906 7783 5962 7792
rect 5540 7754 5592 7760
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5448 5704 5500 5710
rect 5446 5672 5448 5681
rect 5500 5672 5502 5681
rect 5446 5607 5502 5616
rect 5552 3738 5580 7754
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7342 5764 7686
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5906 7304 5962 7313
rect 5906 7239 5962 7248
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 5644 6458 5672 6695
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 5846 5764 6598
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5828 5234 5856 6938
rect 5920 6458 5948 7239
rect 6012 6798 6040 8570
rect 6288 8566 6316 8735
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6104 7857 6132 8434
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6090 7848 6146 7857
rect 6090 7783 6146 7792
rect 6104 7342 6132 7783
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5828 4554 5856 5170
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 6012 4146 6040 6054
rect 6104 4690 6132 7278
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6196 4622 6224 7958
rect 6380 7750 6408 8366
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7472 6328 7478
rect 6380 7449 6408 7686
rect 6276 7414 6328 7420
rect 6366 7440 6422 7449
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 6288 3097 6316 7414
rect 6366 7375 6422 7384
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6380 5642 6408 6870
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6380 4146 6408 4218
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6472 3738 6500 12038
rect 6564 11937 6592 12158
rect 6550 11928 6606 11937
rect 6656 11898 6684 12310
rect 6748 12102 6776 13126
rect 6840 12986 6868 13398
rect 7392 13326 7420 14554
rect 7484 14482 7512 16662
rect 7760 16522 7788 17138
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7838 15464 7894 15473
rect 8036 15434 8064 15506
rect 7838 15399 7840 15408
rect 7892 15399 7894 15408
rect 8024 15428 8076 15434
rect 7840 15370 7892 15376
rect 8024 15370 8076 15376
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7760 14278 7788 14554
rect 8128 14482 8156 16118
rect 8220 15706 8248 16186
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8114 14376 8170 14385
rect 8114 14311 8116 14320
rect 8168 14311 8170 14320
rect 8116 14282 8168 14288
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 7562 13968 7618 13977
rect 7562 13903 7618 13912
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13320 7432 13326
rect 7300 13280 7380 13308
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6932 12628 6960 13126
rect 6840 12600 6960 12628
rect 6736 12096 6788 12102
rect 6840 12073 6868 12600
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6736 12038 6788 12044
rect 6826 12064 6882 12073
rect 6826 11999 6882 12008
rect 6550 11863 6606 11872
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6564 6866 6592 11562
rect 6656 11286 6684 11834
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 11354 6776 11766
rect 6932 11642 6960 12106
rect 6840 11614 6960 11642
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6656 6322 6684 10950
rect 6748 9450 6776 11086
rect 6840 9625 6868 11614
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7208 10606 7236 11222
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6826 9616 6882 9625
rect 6826 9551 6882 9560
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 7024 9382 7052 9658
rect 7300 9586 7328 13280
rect 7380 13262 7432 13268
rect 7484 12306 7512 13806
rect 7576 13190 7604 13903
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7760 12714 7788 12854
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 12442 7604 12582
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 9704 7420 12038
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7470 11928 7526 11937
rect 7610 11931 7918 11940
rect 7564 11892 7616 11898
rect 7526 11872 7564 11880
rect 7470 11863 7564 11872
rect 7484 11852 7564 11863
rect 7564 11834 7616 11840
rect 7746 11792 7802 11801
rect 7746 11727 7802 11736
rect 7930 11792 7986 11801
rect 7930 11727 7986 11736
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7484 9704 7512 11630
rect 7760 11529 7788 11727
rect 7746 11520 7802 11529
rect 7746 11455 7802 11464
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7760 11014 7788 11183
rect 7944 11150 7972 11727
rect 8036 11354 8064 12378
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7932 11144 7984 11150
rect 8128 11098 8156 13330
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8220 12170 8248 13194
rect 8312 12374 8340 16458
rect 8496 16017 8524 17206
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8482 16008 8538 16017
rect 8482 15943 8538 15952
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8404 14414 8432 14758
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8298 12200 8354 12209
rect 8208 12164 8260 12170
rect 8298 12135 8354 12144
rect 8208 12106 8260 12112
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7932 11086 7984 11092
rect 8036 11070 8156 11098
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7944 10606 7972 10746
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 8036 10130 8064 11070
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10674 8156 10950
rect 8220 10810 8248 11834
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8116 10668 8168 10674
rect 8312 10656 8340 12135
rect 8404 11762 8432 14350
rect 8496 12288 8524 15302
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8588 12481 8616 12854
rect 8574 12472 8630 12481
rect 8574 12407 8630 12416
rect 8496 12260 8616 12288
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8116 10610 8168 10616
rect 8220 10628 8340 10656
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 7392 9676 7430 9704
rect 7484 9676 7696 9704
rect 7402 9602 7430 9676
rect 7668 9602 7696 9676
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7392 9574 7430 9602
rect 7484 9574 7696 9602
rect 7748 9580 7800 9586
rect 7012 9376 7064 9382
rect 7116 9364 7144 9522
rect 7392 9364 7420 9574
rect 7116 9336 7328 9364
rect 7392 9336 7430 9364
rect 7012 9318 7064 9324
rect 7300 9330 7328 9336
rect 7300 9302 7334 9330
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 7306 9178 7334 9302
rect 7402 9194 7430 9336
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7392 9166 7430 9194
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6748 4146 6776 8842
rect 6840 8498 6868 8910
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7116 8430 7144 8774
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6932 8276 6960 8366
rect 6840 8248 6960 8276
rect 6840 7936 6868 8248
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 6840 7908 7052 7936
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 7546 6868 7754
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7392 6960 7686
rect 6840 7364 6960 7392
rect 6840 6118 6868 7364
rect 7024 7206 7052 7908
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7116 7274 7144 7346
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6390 7052 6598
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5030 6868 6054
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 7300 4826 7328 8842
rect 7392 6798 7420 9166
rect 7484 7546 7512 9574
rect 7748 9522 7800 9528
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9110 7604 9454
rect 7760 9353 7788 9522
rect 7840 9376 7892 9382
rect 7746 9344 7802 9353
rect 7840 9318 7892 9324
rect 7746 9279 7802 9288
rect 7852 9110 7880 9318
rect 7930 9208 7986 9217
rect 8128 9194 8156 10610
rect 8220 9994 8248 10628
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8496 9722 8524 12106
rect 8588 10656 8616 12260
rect 8680 12102 8708 14010
rect 8772 12102 8800 15642
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8666 11928 8722 11937
rect 8666 11863 8668 11872
rect 8720 11863 8722 11872
rect 8668 11834 8720 11840
rect 8680 11014 8708 11834
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8588 10628 8708 10656
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8588 10441 8616 10474
rect 8680 10470 8708 10628
rect 8668 10464 8720 10470
rect 8574 10432 8630 10441
rect 8668 10406 8720 10412
rect 8574 10367 8630 10376
rect 8680 10305 8708 10406
rect 8666 10296 8722 10305
rect 8666 10231 8722 10240
rect 8666 10024 8722 10033
rect 8576 9988 8628 9994
rect 8666 9959 8668 9968
rect 8576 9930 8628 9936
rect 8720 9959 8722 9968
rect 8668 9930 8720 9936
rect 8588 9761 8616 9930
rect 8574 9752 8630 9761
rect 8484 9716 8536 9722
rect 8574 9687 8630 9696
rect 8484 9658 8536 9664
rect 8220 9450 8432 9466
rect 8208 9444 8432 9450
rect 8260 9438 8432 9444
rect 8208 9386 8260 9392
rect 8404 9382 8432 9438
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7930 9143 7986 9152
rect 8036 9166 8156 9194
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7656 8968 7708 8974
rect 7944 8956 7972 9143
rect 8036 8974 8064 9166
rect 8116 9104 8168 9110
rect 8168 9064 8248 9092
rect 8116 9046 8168 9052
rect 7708 8928 7972 8956
rect 7656 8910 7708 8916
rect 7944 8820 7972 8928
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7944 8792 8064 8820
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 8036 8514 8064 8792
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7944 8486 8064 8514
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 7562 8120 7618 8129
rect 7562 8055 7618 8064
rect 7576 7857 7604 8055
rect 7668 7886 7696 8434
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 7880 7708 7886
rect 7562 7848 7618 7857
rect 7656 7822 7708 7828
rect 7562 7783 7618 7792
rect 7760 7750 7788 8366
rect 7944 8362 7972 8486
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7852 7857 7880 8298
rect 7838 7848 7894 7857
rect 7838 7783 7894 7792
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 7206 7880 7346
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7484 6662 7512 7142
rect 7852 7002 7880 7142
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7654 6352 7710 6361
rect 7654 6287 7710 6296
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7392 5370 7420 5850
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7484 5216 7512 6122
rect 7668 5953 7696 6287
rect 7654 5944 7710 5953
rect 7654 5879 7710 5888
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 8036 5234 8064 8366
rect 8128 7954 8156 8502
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7564 5228 7616 5234
rect 7484 5188 7564 5216
rect 7564 5170 7616 5176
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6840 4622 6868 4762
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 7392 4282 7420 4694
rect 7484 4622 7512 4927
rect 7576 4826 7604 5170
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6274 3088 6330 3097
rect 6274 3023 6330 3032
rect 6840 2854 6868 3878
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 8036 3602 8064 5170
rect 8128 3942 8156 7686
rect 8220 5386 8248 9064
rect 8668 8968 8720 8974
rect 8574 8936 8630 8945
rect 8668 8910 8720 8916
rect 8574 8871 8630 8880
rect 8482 8800 8538 8809
rect 8482 8735 8538 8744
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 5642 8340 7822
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8220 5358 8340 5386
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8220 4010 8248 5238
rect 8312 4690 8340 5358
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8300 4208 8352 4214
rect 8298 4176 8300 4185
rect 8352 4176 8354 4185
rect 8298 4111 8354 4120
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8404 2854 8432 8298
rect 8496 4826 8524 8735
rect 8588 7002 8616 8871
rect 8680 8838 8708 8910
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8673 8708 8774
rect 8666 8664 8722 8673
rect 8666 8599 8722 8608
rect 8666 8256 8722 8265
rect 8666 8191 8722 8200
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8588 6662 8616 6938
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8496 4282 8524 4762
rect 8588 4758 8616 6598
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8680 4282 8708 8191
rect 8772 7954 8800 11630
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8864 6254 8892 12718
rect 8956 9654 8984 13806
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6254 8984 6666
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 9048 5302 9076 13194
rect 9140 10674 9168 14758
rect 9232 12442 9260 16526
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9600 15434 9628 15574
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9312 15088 9364 15094
rect 9310 15056 9312 15065
rect 9416 15076 9444 15302
rect 9496 15088 9548 15094
rect 9364 15056 9366 15065
rect 9310 14991 9366 15000
rect 9416 15048 9496 15076
rect 9416 14618 9444 15048
rect 9496 15030 9548 15036
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11150 9260 12038
rect 9324 11257 9352 12650
rect 9416 11898 9444 13942
rect 9508 11937 9536 14758
rect 9692 13734 9720 17206
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9494 11928 9550 11937
rect 9404 11892 9456 11898
rect 9494 11863 9550 11872
rect 9404 11834 9456 11840
rect 9310 11248 9366 11257
rect 9310 11183 9366 11192
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9140 9110 9168 10066
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9232 8945 9260 11086
rect 9402 10976 9458 10985
rect 9402 10911 9458 10920
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 9126 8392 9182 8401
rect 9232 8362 9260 8871
rect 9324 8838 9352 10610
rect 9416 9654 9444 10911
rect 9508 10742 9536 11154
rect 9600 10849 9628 12582
rect 9678 11248 9734 11257
rect 9678 11183 9734 11192
rect 9692 11082 9720 11183
rect 9784 11082 9812 17274
rect 10416 15632 10468 15638
rect 10322 15600 10378 15609
rect 10416 15574 10468 15580
rect 10322 15535 10378 15544
rect 10336 15502 10364 15535
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10152 13734 10180 15030
rect 10324 14952 10376 14958
rect 10428 14929 10456 15574
rect 10324 14894 10376 14900
rect 10414 14920 10470 14929
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9956 13320 10008 13326
rect 9954 13288 9956 13297
rect 10008 13288 10010 13297
rect 9954 13223 10010 13232
rect 10046 13016 10102 13025
rect 10046 12951 10048 12960
rect 10100 12951 10102 12960
rect 10048 12922 10100 12928
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9876 11642 9904 12378
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9954 11928 10010 11937
rect 9954 11863 10010 11872
rect 9968 11762 9996 11863
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9876 11614 9996 11642
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9586 10840 9642 10849
rect 9586 10775 9642 10784
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9784 10248 9812 11018
rect 9692 10220 9812 10248
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9494 9752 9550 9761
rect 9494 9687 9550 9696
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9353 9444 9454
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 9508 9042 9536 9687
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9126 8327 9182 8336
rect 9220 8356 9272 8362
rect 9140 6798 9168 8327
rect 9220 8298 9272 8304
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9232 5658 9260 8298
rect 9324 6866 9352 8774
rect 9416 8498 9444 8842
rect 9600 8634 9628 9823
rect 9692 9042 9720 10220
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9784 9042 9812 9590
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9508 8362 9536 8570
rect 9692 8430 9720 8978
rect 9680 8424 9732 8430
rect 9678 8392 9680 8401
rect 9732 8392 9734 8401
rect 9496 8356 9548 8362
rect 9678 8327 9734 8336
rect 9496 8298 9548 8304
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 8129 9720 8230
rect 9678 8120 9734 8129
rect 9678 8055 9734 8064
rect 9494 7984 9550 7993
rect 9494 7919 9550 7928
rect 9588 7948 9640 7954
rect 9508 7002 9536 7919
rect 9588 7890 9640 7896
rect 9600 7002 9628 7890
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6730 9536 6802
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9508 5778 9536 6666
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9232 5630 9352 5658
rect 9324 5370 9352 5630
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9324 5098 9352 5306
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9508 5001 9536 5714
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9600 5370 9628 5578
rect 9692 5545 9720 6326
rect 9784 5914 9812 8978
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9494 4992 9550 5001
rect 9494 4927 9550 4936
rect 9600 4622 9628 5306
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 9692 4214 9720 5199
rect 8944 4208 8996 4214
rect 9036 4208 9088 4214
rect 8944 4150 8996 4156
rect 9034 4176 9036 4185
rect 9680 4208 9732 4214
rect 9088 4176 9090 4185
rect 8956 3466 8984 4150
rect 9034 4111 9090 4120
rect 9402 4176 9458 4185
rect 9680 4150 9732 4156
rect 9402 4111 9458 4120
rect 9034 4040 9090 4049
rect 9034 3975 9090 3984
rect 9048 3466 9076 3975
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8680 3058 8708 3402
rect 8956 3126 8984 3402
rect 9232 3210 9260 3538
rect 9310 3496 9366 3505
rect 9310 3431 9366 3440
rect 9324 3398 9352 3431
rect 9416 3398 9444 4111
rect 9588 4072 9640 4078
rect 9508 4020 9588 4026
rect 9508 4014 9640 4020
rect 9508 3998 9628 4014
rect 9508 3670 9536 3998
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9600 3602 9628 3878
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9496 3528 9548 3534
rect 9784 3482 9812 5646
rect 9876 3602 9904 11494
rect 9968 8362 9996 11614
rect 10060 9586 10088 12038
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 8838 10088 9522
rect 10152 9042 10180 13670
rect 10336 13394 10364 14894
rect 10414 14855 10470 14864
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10230 13152 10286 13161
rect 10230 13087 10286 13096
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10138 8800 10194 8809
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9968 7954 9996 8298
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 5302 9996 7890
rect 10060 5710 10088 8774
rect 10138 8735 10194 8744
rect 10152 8312 10180 8735
rect 10244 8362 10272 13087
rect 10336 12782 10364 13330
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12442 10364 12718
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 10130 10364 12106
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10232 8356 10284 8362
rect 10140 8306 10192 8312
rect 10232 8298 10284 8304
rect 10140 8248 10192 8254
rect 10230 8256 10286 8265
rect 10230 8191 10286 8200
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10152 5098 10180 7822
rect 10244 6458 10272 8191
rect 10336 7546 10364 9862
rect 10428 9178 10456 13806
rect 10520 11762 10548 17274
rect 15672 17270 15700 17546
rect 18510 17504 18566 17513
rect 17610 17436 17918 17445
rect 18510 17439 18566 17448
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 18524 17338 18552 17439
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10612 15366 10640 17138
rect 11612 17128 11664 17134
rect 11610 17096 11612 17105
rect 11704 17128 11756 17134
rect 11664 17096 11666 17105
rect 10876 17060 10928 17066
rect 11704 17070 11756 17076
rect 11610 17031 11666 17040
rect 10876 17002 10928 17008
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10598 15056 10654 15065
rect 10598 14991 10654 15000
rect 10612 14958 10640 14991
rect 10600 14952 10652 14958
rect 10704 14940 10732 16186
rect 10888 15065 10916 17002
rect 11716 16998 11744 17070
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11256 15706 11284 15982
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10874 15056 10930 15065
rect 10874 14991 10930 15000
rect 10652 14912 10732 14940
rect 10600 14894 10652 14900
rect 10704 14822 10732 14912
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10612 14521 10640 14758
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10598 13832 10654 13841
rect 10598 13767 10654 13776
rect 10612 12238 10640 13767
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10598 11928 10654 11937
rect 10598 11863 10654 11872
rect 10612 11830 10640 11863
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10520 11354 10548 11494
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 11121 10548 11154
rect 10506 11112 10562 11121
rect 10506 11047 10562 11056
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10810 10548 10950
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10612 10062 10640 11630
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8945 10456 8978
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10414 8800 10470 8809
rect 10414 8735 10470 8744
rect 10428 8566 10456 8735
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 7886 10456 8298
rect 10520 7886 10548 9114
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10612 7698 10640 9998
rect 10704 9926 10732 14758
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 11558 10824 12786
rect 10888 12238 10916 14894
rect 10968 12912 11020 12918
rect 10966 12880 10968 12889
rect 11020 12880 11022 12889
rect 10966 12815 11022 12824
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11072 12170 11100 15506
rect 11256 15502 11284 15642
rect 11716 15502 11744 16594
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11244 15496 11296 15502
rect 11704 15496 11756 15502
rect 11296 15456 11376 15484
rect 11244 15438 11296 15444
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11150 13016 11206 13025
rect 11150 12951 11206 12960
rect 11164 12646 11192 12951
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10888 11558 10916 11698
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11370 10916 11494
rect 10796 11342 10916 11370
rect 10796 9926 10824 11342
rect 11072 11286 11100 12106
rect 11256 11880 11284 14282
rect 11348 14278 11376 15456
rect 11704 15438 11756 15444
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 12050 11376 14214
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11440 12238 11468 13942
rect 11808 13705 11836 16390
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11992 14074 12020 14418
rect 12084 14113 12112 14418
rect 12070 14104 12126 14113
rect 11980 14068 12032 14074
rect 12070 14039 12126 14048
rect 11980 14010 12032 14016
rect 12360 14006 12388 14758
rect 12452 14521 12480 16526
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12438 14512 12494 14521
rect 12438 14447 12494 14456
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12360 13734 12388 13942
rect 12348 13728 12400 13734
rect 11794 13696 11850 13705
rect 12348 13670 12400 13676
rect 11794 13631 11850 13640
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11348 12022 11468 12050
rect 11256 11852 11376 11880
rect 11348 11626 11376 11852
rect 11152 11620 11204 11626
rect 11336 11620 11388 11626
rect 11204 11580 11284 11608
rect 11152 11562 11204 11568
rect 11150 11384 11206 11393
rect 11150 11319 11206 11328
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 11014 11100 11222
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10690 9208 10746 9217
rect 10690 9143 10746 9152
rect 10704 9110 10732 9143
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8809 10732 8842
rect 10690 8800 10746 8809
rect 10690 8735 10746 8744
rect 10428 7670 10640 7698
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10336 7410 10364 7482
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10230 6080 10286 6089
rect 10230 6015 10286 6024
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4622 9996 4966
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9548 3476 9812 3482
rect 9496 3470 9812 3476
rect 9508 3454 9812 3470
rect 9968 3466 9996 3538
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9232 3182 9536 3210
rect 10060 3194 10088 4150
rect 10244 3942 10272 6015
rect 10336 5681 10364 7346
rect 10322 5672 10378 5681
rect 10322 5607 10378 5616
rect 10336 5234 10364 5607
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10336 4826 10364 5034
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10428 4758 10456 7670
rect 10704 7528 10732 8735
rect 10796 8634 10824 9590
rect 10888 8922 10916 10066
rect 10980 9761 11008 10066
rect 10966 9752 11022 9761
rect 10966 9687 11022 9696
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9058 11008 9318
rect 11072 9178 11100 10474
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10980 9030 11100 9058
rect 10888 8894 11008 8922
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10888 8362 10916 8502
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10612 7500 10732 7528
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10520 6497 10548 7414
rect 10612 6934 10640 7500
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 6934 10732 7346
rect 10796 7342 10824 7686
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10506 6488 10562 6497
rect 10506 6423 10562 6432
rect 10612 6254 10640 6598
rect 10690 6488 10746 6497
rect 10690 6423 10746 6432
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10520 5574 10548 6190
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 5552 2446 5580 2790
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 5998 2680 6054 2689
rect 6950 2683 7258 2692
rect 5998 2615 6000 2624
rect 6052 2615 6054 2624
rect 6000 2586 6052 2592
rect 9508 2514 9536 3182
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10520 3126 10548 5510
rect 10612 4826 10640 5578
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10704 4758 10732 6423
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10796 5914 10824 6258
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5846 10916 7822
rect 10980 7478 11008 8894
rect 11072 8294 11100 9030
rect 11164 8945 11192 11319
rect 11256 11082 11284 11580
rect 11336 11562 11388 11568
rect 11334 11520 11390 11529
rect 11334 11455 11390 11464
rect 11348 11082 11376 11455
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11242 10976 11298 10985
rect 11242 10911 11298 10920
rect 11256 9625 11284 10911
rect 11334 10840 11390 10849
rect 11334 10775 11336 10784
rect 11388 10775 11390 10784
rect 11336 10746 11388 10752
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8378 11192 8774
rect 11256 8537 11284 9551
rect 11242 8528 11298 8537
rect 11242 8463 11298 8472
rect 11242 8392 11298 8401
rect 11164 8350 11242 8378
rect 11242 8327 11298 8336
rect 11072 8266 11192 8294
rect 11060 8016 11112 8022
rect 11058 7984 11060 7993
rect 11112 7984 11114 7993
rect 11058 7919 11114 7928
rect 11058 7848 11114 7857
rect 11058 7783 11114 7792
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 6934 11008 7414
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10980 6066 11008 6870
rect 11072 6322 11100 7783
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10980 6038 11100 6066
rect 11072 5953 11100 6038
rect 11058 5944 11114 5953
rect 11058 5879 11114 5888
rect 10876 5840 10928 5846
rect 10782 5808 10838 5817
rect 10876 5782 10928 5788
rect 10782 5743 10838 5752
rect 10796 5642 10824 5743
rect 10966 5672 11022 5681
rect 10784 5636 10836 5642
rect 10966 5607 11022 5616
rect 10784 5578 10836 5584
rect 10980 5574 11008 5607
rect 10968 5568 11020 5574
rect 10782 5536 10838 5545
rect 10968 5510 11020 5516
rect 10782 5471 10838 5480
rect 10796 5370 10824 5471
rect 10874 5400 10930 5409
rect 10784 5364 10836 5370
rect 10874 5335 10930 5344
rect 10784 5306 10836 5312
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10888 4486 10916 5335
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 3194 10916 4422
rect 11072 4282 11100 5879
rect 11164 4758 11192 8266
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 4214 11192 4490
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11256 4078 11284 8327
rect 11348 7449 11376 10746
rect 11440 8906 11468 12022
rect 11532 11354 11560 12922
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12442 11744 12786
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 12256 12640 12308 12646
rect 12360 12628 12388 13670
rect 12452 12850 12480 14350
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12308 12600 12388 12628
rect 12256 12582 12308 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11506 11744 12174
rect 11808 11694 11836 12582
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11624 11478 11744 11506
rect 11796 11552 11848 11558
rect 11900 11540 11928 12378
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11978 11928 12034 11937
rect 11978 11863 11980 11872
rect 12032 11863 12034 11872
rect 11980 11834 12032 11840
rect 12084 11744 12112 12038
rect 12176 11898 12204 12310
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 12050 12296 12242
rect 12440 12096 12492 12102
rect 12268 12022 12388 12050
rect 12440 12038 12492 12044
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12164 11756 12216 11762
rect 12084 11716 12164 11744
rect 12164 11698 12216 11704
rect 11848 11512 11928 11540
rect 11796 11494 11848 11500
rect 11624 11354 11652 11478
rect 11702 11384 11758 11393
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11612 11348 11664 11354
rect 11702 11319 11704 11328
rect 11612 11290 11664 11296
rect 11756 11319 11758 11328
rect 11704 11290 11756 11296
rect 11532 10849 11560 11290
rect 11716 11234 11744 11290
rect 11624 11206 11744 11234
rect 11518 10840 11574 10849
rect 11518 10775 11574 10784
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11532 10577 11560 10678
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11532 9994 11560 10503
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11426 8664 11482 8673
rect 11426 8599 11428 8608
rect 11480 8599 11482 8608
rect 11428 8570 11480 8576
rect 11334 7440 11390 7449
rect 11334 7375 11390 7384
rect 11336 7200 11388 7206
rect 11334 7168 11336 7177
rect 11388 7168 11390 7177
rect 11334 7103 11390 7112
rect 11348 6798 11376 7103
rect 11440 6984 11468 8570
rect 11532 7698 11560 9930
rect 11624 8673 11652 11206
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11610 8664 11666 8673
rect 11610 8599 11666 8608
rect 11610 8120 11666 8129
rect 11610 8055 11612 8064
rect 11664 8055 11666 8064
rect 11612 8026 11664 8032
rect 11532 7670 11652 7698
rect 11518 7576 11574 7585
rect 11518 7511 11574 7520
rect 11532 7478 11560 7511
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11440 6956 11560 6984
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11336 6792 11388 6798
rect 11440 6769 11468 6802
rect 11336 6734 11388 6740
rect 11426 6760 11482 6769
rect 11426 6695 11482 6704
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 6118 11376 6598
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 4072 11296 4078
rect 10966 4040 11022 4049
rect 11244 4014 11296 4020
rect 10966 3975 11022 3984
rect 10980 3534 11008 3975
rect 11348 3670 11376 5102
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 10968 3528 11020 3534
rect 11532 3482 11560 6956
rect 11624 6100 11652 7670
rect 11716 6662 11744 11086
rect 11808 10198 11836 11494
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12176 10452 12204 11290
rect 12360 11014 12388 12022
rect 12452 11762 12480 12038
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12348 11008 12400 11014
rect 12452 10985 12480 11562
rect 12348 10950 12400 10956
rect 12438 10976 12494 10985
rect 12268 10606 12296 10950
rect 12438 10911 12494 10920
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12452 10742 12480 10775
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12176 10424 12388 10452
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 12360 10130 12388 10424
rect 12438 10160 12494 10169
rect 12348 10124 12400 10130
rect 12438 10095 12494 10104
rect 12348 10066 12400 10072
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12346 9888 12402 9897
rect 11796 9512 11848 9518
rect 12268 9489 12296 9862
rect 12346 9823 12402 9832
rect 11796 9454 11848 9460
rect 12254 9480 12310 9489
rect 11808 9042 11836 9454
rect 12254 9415 12310 9424
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 7954 11836 8978
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8430 11928 8842
rect 11992 8809 12020 9114
rect 12360 9092 12388 9823
rect 12176 9064 12388 9092
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 12176 8566 12204 9064
rect 12254 8936 12310 8945
rect 12254 8871 12256 8880
rect 12308 8871 12310 8880
rect 12256 8842 12308 8848
rect 12346 8800 12402 8809
rect 12346 8735 12402 8744
rect 12360 8566 12388 8735
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7721 11836 7890
rect 11888 7744 11940 7750
rect 11794 7712 11850 7721
rect 11888 7686 11940 7692
rect 12452 7698 12480 10095
rect 12544 8378 12572 16458
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15638 12664 15846
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12728 13569 12756 13738
rect 12714 13560 12770 13569
rect 12714 13495 12770 13504
rect 12820 13190 12848 13738
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13530 12940 13670
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12636 12170 12664 12310
rect 12808 12232 12860 12238
rect 12806 12200 12808 12209
rect 12860 12200 12862 12209
rect 12624 12164 12676 12170
rect 12806 12135 12862 12144
rect 12912 12152 12940 12786
rect 13004 12220 13032 15982
rect 13188 15706 13216 16594
rect 13280 16114 13308 16934
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13082 15600 13138 15609
rect 13082 15535 13138 15544
rect 13096 12288 13124 15535
rect 13280 14006 13308 16050
rect 13372 15638 13400 16390
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13096 12260 13216 12288
rect 13004 12192 13124 12220
rect 12912 12124 13032 12152
rect 12624 12106 12676 12112
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12636 11218 12664 11834
rect 13004 11762 13032 12124
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12728 11354 12756 11698
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 13004 10577 13032 11698
rect 13096 11014 13124 12192
rect 13188 12102 13216 12260
rect 13280 12238 13308 13738
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12990 10568 13046 10577
rect 12990 10503 13046 10512
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12636 9586 12664 9658
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 13004 8634 13032 9658
rect 13096 9586 13124 10406
rect 13188 9586 13216 11154
rect 13280 10674 13308 11630
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13096 9466 13124 9522
rect 13096 9438 13308 9466
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13082 8528 13138 8537
rect 12992 8492 13044 8498
rect 13082 8463 13138 8472
rect 12992 8434 13044 8440
rect 12544 8350 12756 8378
rect 12728 7818 12756 8350
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12912 7750 12940 8026
rect 12900 7744 12952 7750
rect 11794 7647 11850 7656
rect 11808 7546 11836 7647
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11900 7188 11928 7686
rect 12452 7670 12572 7698
rect 12900 7686 12952 7692
rect 11808 7160 11928 7188
rect 12348 7200 12400 7206
rect 11808 6780 11836 7160
rect 12348 7142 12400 7148
rect 12544 7154 12572 7670
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12622 7168 12678 7177
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11888 6792 11940 6798
rect 11808 6752 11888 6780
rect 12072 6792 12124 6798
rect 11888 6734 11940 6740
rect 11992 6740 12072 6746
rect 11992 6734 12124 6740
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11702 6488 11758 6497
rect 11900 6458 11928 6734
rect 11992 6718 12112 6734
rect 11992 6662 12020 6718
rect 12176 6662 12204 6938
rect 12360 6866 12388 7142
rect 12544 7126 12622 7154
rect 12622 7103 12678 7112
rect 12636 7002 12664 7103
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 11702 6423 11758 6432
rect 11888 6452 11940 6458
rect 11716 6390 11744 6423
rect 11888 6394 11940 6400
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11704 6248 11756 6254
rect 11756 6196 12204 6202
rect 11704 6190 12204 6196
rect 11716 6186 12204 6190
rect 11716 6180 12216 6186
rect 11716 6174 12164 6180
rect 12164 6122 12216 6128
rect 12268 6118 12296 6666
rect 12452 6633 12480 6734
rect 12438 6624 12494 6633
rect 12438 6559 12494 6568
rect 12544 6440 12572 6938
rect 12820 6662 12848 7210
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 13004 6440 13032 8434
rect 13096 8430 13124 8463
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12544 6412 12664 6440
rect 12636 6186 12664 6412
rect 12820 6412 13032 6440
rect 12714 6352 12770 6361
rect 12714 6287 12770 6296
rect 12728 6186 12756 6287
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12072 6112 12124 6118
rect 11624 6072 12072 6100
rect 12072 6054 12124 6060
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 12544 5914 12572 6054
rect 12532 5908 12584 5914
rect 12584 5868 12664 5896
rect 12532 5850 12584 5856
rect 12530 5808 12586 5817
rect 12636 5778 12664 5868
rect 12530 5743 12586 5752
rect 12624 5772 12676 5778
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11624 4214 11652 5238
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11702 3768 11758 3777
rect 11702 3703 11758 3712
rect 11716 3534 11744 3703
rect 11808 3618 11836 4014
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11808 3590 11928 3618
rect 11900 3534 11928 3590
rect 10968 3470 11020 3476
rect 11440 3454 11560 3482
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10888 3058 10916 3130
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11440 2650 11468 3454
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11532 3126 11560 3334
rect 11716 3194 11744 3470
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11716 2582 11744 3130
rect 11808 3058 11836 3470
rect 11900 3058 11928 3470
rect 12084 3126 12112 3674
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 11808 2310 11836 2994
rect 11900 2922 11928 2994
rect 12176 2922 12204 3334
rect 12544 3210 12572 5743
rect 12624 5714 12676 5720
rect 12820 5642 12848 6412
rect 13096 6372 13124 8366
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13004 6344 13124 6372
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12912 5953 12940 6258
rect 12898 5944 12954 5953
rect 12898 5879 12954 5888
rect 12898 5808 12954 5817
rect 12898 5743 12954 5752
rect 12912 5710 12940 5743
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13004 4706 13032 6344
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13096 5914 13124 6122
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 13096 5370 13124 5578
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4826 13124 4966
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13004 4678 13124 4706
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12990 4176 13046 4185
rect 12990 4111 12992 4120
rect 13044 4111 13046 4120
rect 12992 4082 13044 4088
rect 12992 3392 13044 3398
rect 13096 3380 13124 4678
rect 13044 3352 13124 3380
rect 12992 3334 13044 3340
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 12452 3182 12572 3210
rect 12452 3126 12480 3182
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 13004 3058 13032 3334
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 13188 2378 13216 8298
rect 13280 6202 13308 9438
rect 13372 8634 13400 14554
rect 13464 12345 13492 17206
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 13740 17105 13768 17138
rect 13726 17096 13782 17105
rect 13726 17031 13782 17040
rect 14384 16998 14412 17138
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13556 13938 13584 14418
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13648 13818 13676 15370
rect 14016 15162 14044 16730
rect 14186 16688 14242 16697
rect 14186 16623 14188 16632
rect 14240 16623 14242 16632
rect 14188 16594 14240 16600
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 13556 13790 13676 13818
rect 13450 12336 13506 12345
rect 13450 12271 13506 12280
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 12102 13492 12174
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 9110 13492 12038
rect 13556 11286 13584 13790
rect 13740 13394 13768 15098
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13832 13326 13860 13874
rect 13924 13433 13952 14758
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 13910 13424 13966 13433
rect 13910 13359 13966 13368
rect 13820 13320 13872 13326
rect 13634 13288 13690 13297
rect 13820 13262 13872 13268
rect 13634 13223 13636 13232
rect 13688 13223 13690 13232
rect 13636 13194 13688 13200
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13634 12064 13690 12073
rect 13634 11999 13690 12008
rect 13648 11830 13676 11999
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13372 7410 13400 8026
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13372 7018 13400 7346
rect 13464 7206 13492 8298
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13372 6990 13492 7018
rect 13464 6304 13492 6990
rect 13556 6372 13584 11086
rect 13648 7732 13676 11222
rect 13740 8090 13768 12786
rect 13832 12170 13860 13262
rect 14108 13161 14136 13942
rect 14094 13152 14150 13161
rect 14094 13087 14150 13096
rect 13910 12744 13966 12753
rect 13910 12679 13912 12688
rect 13964 12679 13966 12688
rect 13912 12650 13964 12656
rect 13910 12608 13966 12617
rect 13910 12543 13966 12552
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13832 11898 13860 12106
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13818 11112 13874 11121
rect 13818 11047 13820 11056
rect 13872 11047 13874 11056
rect 13820 11018 13872 11024
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 8498 13860 9590
rect 13924 9178 13952 12543
rect 14094 11928 14150 11937
rect 14094 11863 14096 11872
rect 14148 11863 14150 11872
rect 14096 11834 14148 11840
rect 14094 11792 14150 11801
rect 14094 11727 14150 11736
rect 14108 11098 14136 11727
rect 14016 11070 14136 11098
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7857 13768 7890
rect 13726 7848 13782 7857
rect 13726 7783 13782 7792
rect 13648 7704 13768 7732
rect 13634 7576 13690 7585
rect 13634 7511 13690 7520
rect 13648 7478 13676 7511
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6662 13676 7142
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13556 6344 13676 6372
rect 13464 6276 13584 6304
rect 13280 6174 13492 6202
rect 13360 5840 13412 5846
rect 13280 5800 13360 5828
rect 13280 5642 13308 5800
rect 13360 5782 13412 5788
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 5386 13400 5578
rect 13280 5358 13400 5386
rect 13280 5030 13308 5358
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4622 13308 4966
rect 13464 4690 13492 6174
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13556 3942 13584 6276
rect 13648 5846 13676 6344
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13740 4214 13768 7704
rect 13832 7274 13860 8026
rect 13924 7886 13952 8910
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13924 6866 13952 7822
rect 14016 7342 14044 11070
rect 14200 8634 14228 15030
rect 14292 8974 14320 15302
rect 14384 14482 14412 16934
rect 14660 16726 14688 16934
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16114 14872 16458
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14476 15502 14504 15846
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14384 12442 14412 14418
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14384 12238 14412 12378
rect 14372 12232 14424 12238
rect 14370 12200 14372 12209
rect 14424 12200 14426 12209
rect 14370 12135 14426 12144
rect 14370 11928 14426 11937
rect 14370 11863 14426 11872
rect 14384 11286 14412 11863
rect 14476 11694 14504 15438
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 12782 14688 13330
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14752 12434 14780 15846
rect 14844 15094 14872 16050
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14844 14822 14872 15030
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14844 13002 14872 14758
rect 14936 13161 14964 16390
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 13274 15056 15302
rect 15212 15162 15240 16118
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 15042 15332 15506
rect 15212 15014 15332 15042
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15120 13394 15148 14350
rect 15212 13938 15240 15014
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15304 13841 15332 14282
rect 15290 13832 15346 13841
rect 15290 13767 15346 13776
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15292 13320 15344 13326
rect 15028 13246 15148 13274
rect 15292 13262 15344 13268
rect 14922 13152 14978 13161
rect 14922 13087 14978 13096
rect 14844 12974 15056 13002
rect 14922 12880 14978 12889
rect 14922 12815 14978 12824
rect 14660 12406 14780 12434
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 6254 13860 6666
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5642 13860 6054
rect 13924 5710 13952 6394
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5370 13860 5578
rect 13924 5370 13952 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13818 4856 13874 4865
rect 13818 4791 13874 4800
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13832 3670 13860 4791
rect 14016 4282 14044 6938
rect 14108 6458 14136 8570
rect 14292 8498 14320 8774
rect 14384 8634 14412 11086
rect 14476 10470 14504 11086
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14568 9654 14596 12174
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14384 8401 14412 8570
rect 14370 8392 14426 8401
rect 14370 8327 14426 8336
rect 14660 7750 14688 12406
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11354 14872 11494
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 8498 14780 10542
rect 14936 10452 14964 12815
rect 15028 11676 15056 12974
rect 15120 11801 15148 13246
rect 15304 12850 15332 13262
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 15304 11694 15332 12038
rect 15292 11688 15344 11694
rect 15028 11648 15148 11676
rect 14936 10424 15056 10452
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6361 14228 7686
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14278 7032 14334 7041
rect 14278 6967 14334 6976
rect 14292 6390 14320 6967
rect 14384 6730 14412 7210
rect 14648 6928 14700 6934
rect 14554 6896 14610 6905
rect 14648 6870 14700 6876
rect 14554 6831 14556 6840
rect 14608 6831 14610 6840
rect 14556 6802 14608 6808
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14280 6384 14332 6390
rect 14186 6352 14242 6361
rect 14280 6326 14332 6332
rect 14186 6287 14242 6296
rect 14384 5778 14412 6666
rect 14660 6662 14688 6870
rect 14752 6866 14780 8434
rect 14936 7546 14964 10202
rect 15028 8090 15056 10424
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14844 6798 14872 7210
rect 14936 6934 14964 7482
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 14384 3194 14412 5714
rect 14936 4672 14964 6870
rect 15028 6798 15056 7822
rect 15120 7478 15148 11648
rect 15292 11630 15344 11636
rect 15200 11280 15252 11286
rect 15198 11248 15200 11257
rect 15252 11248 15254 11257
rect 15198 11183 15254 11192
rect 15198 9616 15254 9625
rect 15198 9551 15254 9560
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15120 6798 15148 7278
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14844 4644 14964 4672
rect 14844 4078 14872 4644
rect 14922 4584 14978 4593
rect 14922 4519 14924 4528
rect 14976 4519 14978 4528
rect 14924 4490 14976 4496
rect 15028 4486 15056 6734
rect 15212 6458 15240 9551
rect 15304 9042 15332 11630
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15396 8922 15424 15846
rect 15488 12782 15516 16050
rect 15672 15434 15700 16526
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 15094 15608 15302
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15580 12918 15608 15030
rect 15672 13870 15700 15370
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 14006 15792 14418
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13864 15712 13870
rect 15752 13864 15804 13870
rect 15660 13806 15712 13812
rect 15750 13832 15752 13841
rect 15804 13832 15806 13841
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 11150 15516 12718
rect 15672 12434 15700 13806
rect 15750 13767 15806 13776
rect 15856 13002 15884 15642
rect 16028 14884 16080 14890
rect 16028 14826 16080 14832
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15948 13977 15976 14010
rect 15934 13968 15990 13977
rect 15934 13903 15990 13912
rect 16040 13716 16068 14826
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 14074 16252 14214
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16132 13841 16160 13874
rect 16118 13832 16174 13841
rect 16118 13767 16174 13776
rect 16316 13734 16344 15846
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16304 13728 16356 13734
rect 16040 13688 16160 13716
rect 16132 13530 16160 13688
rect 16304 13670 16356 13676
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 15856 12974 16068 13002
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15672 12406 15792 12434
rect 15658 12336 15714 12345
rect 15658 12271 15714 12280
rect 15672 11762 15700 12271
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15488 10742 15516 10950
rect 15476 10736 15528 10742
rect 15580 10713 15608 11562
rect 15672 11393 15700 11562
rect 15658 11384 15714 11393
rect 15658 11319 15714 11328
rect 15476 10678 15528 10684
rect 15566 10704 15622 10713
rect 15566 10639 15622 10648
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15304 8894 15424 8922
rect 15304 8022 15332 8894
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 15304 7546 15332 7958
rect 15382 7576 15438 7585
rect 15292 7540 15344 7546
rect 15382 7511 15438 7520
rect 15292 7482 15344 7488
rect 15396 7478 15424 7511
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15120 5914 15148 6326
rect 15304 6322 15332 7103
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15396 6730 15424 6870
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15304 5914 15332 6258
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15120 4758 15148 5850
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15120 4554 15148 4694
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14384 2378 14412 3130
rect 14924 2576 14976 2582
rect 14922 2544 14924 2553
rect 14976 2544 14978 2553
rect 14922 2479 14978 2488
rect 15120 2446 15148 3130
rect 15212 2650 15240 4762
rect 15304 4758 15332 5850
rect 15488 5030 15516 9522
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 15304 4554 15332 4694
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15580 4282 15608 9046
rect 15672 7274 15700 10610
rect 15764 7886 15792 12406
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 10266 15884 12038
rect 15948 11150 15976 12854
rect 16040 12102 16068 12974
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 11937 16068 12038
rect 16026 11928 16082 11937
rect 16026 11863 16082 11872
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 16040 11014 16068 11630
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 9926 15976 10678
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15672 6440 15700 7210
rect 15764 6798 15792 7822
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15672 6412 15792 6440
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 5778 15700 6258
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15764 5642 15792 6412
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15764 3194 15792 5578
rect 15856 5370 15884 9522
rect 15948 9110 15976 9862
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15948 5234 15976 7210
rect 16040 6798 16068 10950
rect 16132 7274 16160 13466
rect 16316 12918 16344 13670
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16212 12776 16264 12782
rect 16408 12730 16436 14214
rect 16212 12718 16264 12724
rect 16224 12617 16252 12718
rect 16316 12702 16436 12730
rect 16210 12608 16266 12617
rect 16210 12543 16266 12552
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16224 11762 16252 11834
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 10742 16252 11698
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16118 6624 16174 6633
rect 16040 6322 16068 6598
rect 16118 6559 16174 6568
rect 16132 6390 16160 6559
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16040 5001 16068 6258
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5273 16160 6054
rect 16118 5264 16174 5273
rect 16118 5199 16174 5208
rect 16120 5024 16172 5030
rect 16026 4992 16082 5001
rect 16120 4966 16172 4972
rect 16026 4927 16082 4936
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15212 2530 15240 2586
rect 15212 2502 15332 2530
rect 16132 2514 16160 4966
rect 16224 3398 16252 10134
rect 16316 7206 16344 12702
rect 16500 12628 16528 14894
rect 16592 13258 16620 15574
rect 16670 15464 16726 15473
rect 16670 15399 16726 15408
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16580 12912 16632 12918
rect 16684 12889 16712 15399
rect 16580 12854 16632 12860
rect 16670 12880 16726 12889
rect 16408 12600 16528 12628
rect 16408 11898 16436 12600
rect 16592 12434 16620 12854
rect 16670 12815 16726 12824
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16500 12406 16620 12434
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16408 9586 16436 11630
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16394 7440 16450 7449
rect 16394 7375 16450 7384
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16408 3738 16436 7375
rect 16500 5658 16528 12406
rect 16580 12232 16632 12238
rect 16578 12200 16580 12209
rect 16632 12200 16634 12209
rect 16578 12135 16634 12144
rect 16592 11257 16620 12135
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16592 7750 16620 11086
rect 16684 7818 16712 12650
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16592 5778 16620 6326
rect 16684 6322 16712 7754
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16500 5630 16620 5658
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16500 4826 16528 5238
rect 16592 5234 16620 5630
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4826 16620 5034
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16684 4010 16712 6122
rect 16776 5370 16804 16934
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 18512 16448 18564 16454
rect 18510 16416 18512 16425
rect 18564 16416 18566 16425
rect 17610 16348 17918 16357
rect 18510 16351 18566 16360
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17328 14385 17356 14486
rect 17314 14376 17370 14385
rect 16856 14340 16908 14346
rect 17314 14311 17370 14320
rect 16856 14282 16908 14288
rect 16868 12442 16896 14282
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16948 12436 17000 12442
rect 17328 12434 17356 13806
rect 17420 13530 17448 15982
rect 18512 15360 18564 15366
rect 18510 15328 18512 15337
rect 18564 15328 18566 15337
rect 17610 15260 17918 15269
rect 18510 15263 18566 15272
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17512 13376 17540 14418
rect 18236 14272 18288 14278
rect 18234 14240 18236 14249
rect 18288 14240 18290 14249
rect 17610 14172 17918 14181
rect 18234 14175 18290 14184
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 13954 18000 14010
rect 17880 13926 18000 13954
rect 17880 13530 17908 13926
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18156 13530 18184 13806
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 16948 12378 17000 12384
rect 17236 12406 17356 12434
rect 17420 13348 17540 13376
rect 16960 11540 16988 12378
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11937 17080 12038
rect 17038 11928 17094 11937
rect 17038 11863 17094 11872
rect 17236 11694 17264 12406
rect 17316 12096 17368 12102
rect 17314 12064 17316 12073
rect 17368 12064 17370 12073
rect 17314 11999 17370 12008
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16868 11512 16988 11540
rect 16868 9722 16896 11512
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16946 11248 17002 11257
rect 16946 11183 17002 11192
rect 16960 10742 16988 11183
rect 17052 11150 17080 11290
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10810 17080 10950
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16868 6914 16896 9386
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 17328 7834 17356 11766
rect 17420 11082 17448 13348
rect 17604 13172 17632 13466
rect 17512 13144 17632 13172
rect 17512 12442 17540 13144
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12442 17632 12582
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17406 10976 17462 10985
rect 17406 10911 17462 10920
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 17236 7806 17356 7834
rect 16960 7410 16988 7754
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17236 7256 17264 7806
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 7546 17356 7686
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17236 7228 17356 7256
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16868 6886 16988 6914
rect 16960 6322 16988 6886
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 17144 6390 17172 6666
rect 17328 6610 17356 7228
rect 17236 6582 17356 6610
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16854 6216 16910 6225
rect 16854 6151 16856 6160
rect 16908 6151 16910 6160
rect 17236 6168 17264 6582
rect 17314 6488 17370 6497
rect 17314 6423 17316 6432
rect 17368 6423 17370 6432
rect 17316 6394 17368 6400
rect 17420 6390 17448 10911
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17236 6140 17356 6168
rect 16856 6122 16908 6128
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 17144 5166 17172 5578
rect 17236 5370 17264 5850
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 16948 5160 17000 5166
rect 16854 5128 16910 5137
rect 16948 5102 17000 5108
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 16854 5063 16910 5072
rect 16868 4826 16896 5063
rect 16960 5030 16988 5102
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 17328 3466 17356 6140
rect 17420 5914 17448 6326
rect 17512 6322 17540 12242
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17604 11014 17632 11290
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10010 17908 10406
rect 17972 10130 18000 13466
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17880 9982 18000 10010
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17972 9602 18000 9982
rect 17880 9574 18000 9602
rect 17880 8922 17908 9574
rect 17880 8894 18000 8922
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 17972 8548 18000 8894
rect 17880 8520 18000 8548
rect 17880 7732 17908 8520
rect 17880 7704 18000 7732
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 17972 7426 18000 7704
rect 17880 7398 18000 7426
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17604 7002 17632 7142
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17880 6712 17908 7398
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 7002 18000 7210
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18064 6769 18092 12786
rect 18156 12306 18184 13330
rect 18512 13184 18564 13190
rect 18510 13152 18512 13161
rect 18564 13152 18566 13161
rect 18510 13087 18566 13096
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18156 7886 18184 11154
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18050 6760 18106 6769
rect 17880 6684 18000 6712
rect 18050 6695 18106 6704
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17972 6440 18000 6684
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17604 6412 18000 6440
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17604 5794 17632 6412
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17420 5766 17632 5794
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 17420 2922 17448 5766
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 5234 17540 5646
rect 17788 5642 17816 6190
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 18064 5370 18092 6598
rect 18156 6322 18184 6938
rect 18248 6798 18276 12378
rect 18512 12096 18564 12102
rect 18510 12064 18512 12073
rect 18564 12064 18566 12073
rect 18510 11999 18566 12008
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18234 6352 18290 6361
rect 18144 6316 18196 6322
rect 18234 6287 18236 6296
rect 18144 6258 18196 6264
rect 18288 6287 18290 6296
rect 18236 6258 18288 6264
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 18340 4826 18368 11591
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10985 18552 11018
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18432 8945 18460 10066
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18524 9897 18552 9998
rect 18510 9888 18566 9897
rect 18510 9823 18566 9832
rect 18418 8936 18474 8945
rect 18418 8871 18474 8880
rect 18420 8832 18472 8838
rect 18418 8800 18420 8809
rect 18472 8800 18474 8809
rect 18418 8735 18474 8744
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18420 7744 18472 7750
rect 18418 7712 18420 7721
rect 18472 7712 18474 7721
rect 18418 7647 18474 7656
rect 18524 6730 18552 8230
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18420 6656 18472 6662
rect 18418 6624 18420 6633
rect 18472 6624 18474 6633
rect 18418 6559 18474 6568
rect 18420 5568 18472 5574
rect 18418 5536 18420 5545
rect 18472 5536 18474 5545
rect 18418 5471 18474 5480
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18234 4720 18290 4729
rect 18234 4655 18290 4664
rect 18248 4622 18276 4655
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 18156 4214 18184 4490
rect 18420 4480 18472 4486
rect 18418 4448 18420 4457
rect 18472 4448 18474 4457
rect 18418 4383 18474 4392
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 17880 3641 17908 3878
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 18156 3097 18184 3878
rect 18420 3392 18472 3398
rect 18418 3360 18420 3369
rect 18472 3360 18474 3369
rect 18418 3295 18474 3304
rect 18142 3088 18198 3097
rect 18142 3023 18198 3032
rect 17408 2916 17460 2922
rect 17408 2858 17460 2864
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 15304 2446 15332 2502
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 18616 2446 18644 14758
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18786 12744 18842 12753
rect 18786 12679 18842 12688
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18708 4758 18736 8842
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18708 4146 18736 4694
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18800 3534 18828 12679
rect 18892 5681 18920 14350
rect 18878 5672 18934 5681
rect 18878 5607 18934 5616
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 11796 2304 11848 2310
rect 18420 2304 18472 2310
rect 11796 2246 11848 2252
rect 18418 2272 18420 2281
rect 18472 2272 18474 2281
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 17610 2204 17918 2213
rect 18418 2207 18474 2216
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
<< via2 >>
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1582 15036 1584 15056
rect 1584 15036 1636 15056
rect 1636 15036 1638 15056
rect 1582 15000 1638 15036
rect 1398 13368 1454 13424
rect 1582 12688 1638 12744
rect 1674 9560 1730 9616
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 2134 15272 2190 15328
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1950 8372 1952 8392
rect 1952 8372 2004 8392
rect 2004 8372 2006 8392
rect 1950 8336 2006 8372
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3330 16632 3386 16688
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 3146 15136 3202 15192
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2594 13232 2650 13288
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2594 10648 2650 10704
rect 2410 9424 2466 9480
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 3054 12708 3110 12744
rect 3054 12688 3056 12708
rect 3056 12688 3108 12708
rect 3108 12688 3110 12708
rect 3054 9696 3110 9752
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2686 7384 2742 7440
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1398 3984 1454 4040
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3054 7384 3110 7440
rect 3146 6296 3202 6352
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 3514 8200 3570 8256
rect 3514 6996 3570 7032
rect 3514 6976 3516 6996
rect 3516 6976 3568 6996
rect 3568 6976 3570 6996
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3698 12960 3754 13016
rect 4066 13948 4068 13968
rect 4068 13948 4120 13968
rect 4120 13948 4122 13968
rect 4066 13912 4122 13948
rect 3698 11500 3700 11520
rect 3700 11500 3752 11520
rect 3752 11500 3754 11520
rect 3698 11464 3754 11500
rect 3882 7928 3938 7984
rect 3882 7792 3938 7848
rect 4066 10512 4122 10568
rect 4434 13368 4490 13424
rect 4526 11756 4582 11792
rect 4526 11736 4528 11756
rect 4528 11736 4580 11756
rect 4580 11736 4582 11756
rect 4342 10104 4398 10160
rect 4526 9560 4582 9616
rect 4066 8880 4122 8936
rect 4066 8608 4122 8664
rect 4342 9016 4398 9072
rect 4250 8608 4306 8664
rect 4158 8492 4214 8528
rect 4158 8472 4160 8492
rect 4160 8472 4212 8492
rect 4212 8472 4214 8492
rect 4250 8336 4306 8392
rect 4894 15428 4950 15464
rect 4894 15408 4896 15428
rect 4896 15408 4948 15428
rect 4948 15408 4950 15428
rect 5446 15544 5502 15600
rect 4710 12144 4766 12200
rect 4802 8336 4858 8392
rect 4802 6724 4858 6760
rect 4802 6704 4804 6724
rect 4804 6704 4856 6724
rect 4856 6704 4858 6724
rect 5630 13504 5686 13560
rect 5630 11600 5686 11656
rect 5354 8336 5410 8392
rect 5722 8200 5778 8256
rect 6090 15272 6146 15328
rect 5998 9560 6054 9616
rect 5354 6160 5410 6216
rect 5354 6024 5410 6080
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6366 15564 6422 15600
rect 6366 15544 6368 15564
rect 6368 15544 6420 15564
rect 6420 15544 6422 15564
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6734 13776 6790 13832
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 6550 13096 6606 13152
rect 6366 9696 6422 9752
rect 6274 8880 6330 8936
rect 5998 8744 6054 8800
rect 6274 8744 6330 8800
rect 5906 7792 5962 7848
rect 5446 5652 5448 5672
rect 5448 5652 5500 5672
rect 5500 5652 5502 5672
rect 5446 5616 5502 5652
rect 5906 7248 5962 7304
rect 5630 6704 5686 6760
rect 6090 7792 6146 7848
rect 5354 3576 5410 3632
rect 6366 7384 6422 7440
rect 6550 11872 6606 11928
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7838 15428 7894 15464
rect 7838 15408 7840 15428
rect 7840 15408 7892 15428
rect 7892 15408 7894 15428
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 8114 14340 8170 14376
rect 8114 14320 8116 14340
rect 8116 14320 8168 14340
rect 8168 14320 8170 14340
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7562 13912 7618 13968
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6826 12008 6882 12064
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6826 9560 6882 9616
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7470 11872 7526 11928
rect 7746 11736 7802 11792
rect 7930 11736 7986 11792
rect 7746 11464 7802 11520
rect 7746 11192 7802 11248
rect 8482 15952 8538 16008
rect 8298 12144 8354 12200
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 8574 12416 8630 12472
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7746 9288 7802 9344
rect 7930 9152 7986 9208
rect 8666 11892 8722 11928
rect 8666 11872 8668 11892
rect 8668 11872 8720 11892
rect 8720 11872 8722 11892
rect 8574 10376 8630 10432
rect 8666 10240 8722 10296
rect 8666 9988 8722 10024
rect 8666 9968 8668 9988
rect 8668 9968 8720 9988
rect 8720 9968 8722 9988
rect 8574 9696 8630 9752
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7562 8064 7618 8120
rect 7562 7792 7618 7848
rect 7838 7792 7894 7848
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7654 6296 7710 6352
rect 7654 5888 7710 5944
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7470 4936 7526 4992
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6274 3032 6330 3088
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 8574 8880 8630 8936
rect 8482 8744 8538 8800
rect 8298 4156 8300 4176
rect 8300 4156 8352 4176
rect 8352 4156 8354 4176
rect 8298 4120 8354 4156
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 8666 8608 8722 8664
rect 8666 8200 8722 8256
rect 9310 15036 9312 15056
rect 9312 15036 9364 15056
rect 9364 15036 9366 15056
rect 9310 15000 9366 15036
rect 9494 11872 9550 11928
rect 9310 11192 9366 11248
rect 9402 10920 9458 10976
rect 9218 8880 9274 8936
rect 9126 8336 9182 8392
rect 9678 11192 9734 11248
rect 10322 15544 10378 15600
rect 9954 13268 9956 13288
rect 9956 13268 10008 13288
rect 10008 13268 10010 13288
rect 9954 13232 10010 13268
rect 10046 12980 10102 13016
rect 10046 12960 10048 12980
rect 10048 12960 10100 12980
rect 10100 12960 10102 12980
rect 9954 11872 10010 11928
rect 9586 10784 9642 10840
rect 9586 9832 9642 9888
rect 9494 9696 9550 9752
rect 9402 9288 9458 9344
rect 9678 8372 9680 8392
rect 9680 8372 9732 8392
rect 9732 8372 9734 8392
rect 9678 8336 9734 8372
rect 9678 8064 9734 8120
rect 9494 7928 9550 7984
rect 9678 5480 9734 5536
rect 9494 4936 9550 4992
rect 9678 5208 9734 5264
rect 9034 4156 9036 4176
rect 9036 4156 9088 4176
rect 9088 4156 9090 4176
rect 9034 4120 9090 4156
rect 9402 4120 9458 4176
rect 9034 3984 9090 4040
rect 9310 3440 9366 3496
rect 10414 14864 10470 14920
rect 10230 13096 10286 13152
rect 10138 8744 10194 8800
rect 10230 8200 10286 8256
rect 18510 17448 18566 17504
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 11610 17076 11612 17096
rect 11612 17076 11664 17096
rect 11664 17076 11666 17096
rect 11610 17040 11666 17076
rect 10598 15000 10654 15056
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 10874 15000 10930 15056
rect 10598 14456 10654 14512
rect 10598 13776 10654 13832
rect 10598 11872 10654 11928
rect 10506 11056 10562 11112
rect 10414 8880 10470 8936
rect 10414 8744 10470 8800
rect 10966 12860 10968 12880
rect 10968 12860 11020 12880
rect 11020 12860 11022 12880
rect 10966 12824 11022 12860
rect 11150 12960 11206 13016
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 12070 14048 12126 14104
rect 12438 14456 12494 14512
rect 11794 13640 11850 13696
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 11150 11328 11206 11384
rect 10690 9152 10746 9208
rect 10690 8744 10746 8800
rect 10230 6024 10286 6080
rect 10322 5616 10378 5672
rect 10966 9696 11022 9752
rect 10506 6432 10562 6488
rect 10690 6432 10746 6488
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 5998 2644 6054 2680
rect 5998 2624 6000 2644
rect 6000 2624 6052 2644
rect 6052 2624 6054 2644
rect 11334 11464 11390 11520
rect 11242 10920 11298 10976
rect 11334 10804 11390 10840
rect 11334 10784 11336 10804
rect 11336 10784 11388 10804
rect 11388 10784 11390 10804
rect 11242 9560 11298 9616
rect 11150 8880 11206 8936
rect 11242 8472 11298 8528
rect 11242 8336 11298 8392
rect 11058 7964 11060 7984
rect 11060 7964 11112 7984
rect 11112 7964 11114 7984
rect 11058 7928 11114 7964
rect 11058 7792 11114 7848
rect 11058 5888 11114 5944
rect 10782 5752 10838 5808
rect 10966 5616 11022 5672
rect 10782 5480 10838 5536
rect 10874 5344 10930 5400
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11978 11892 12034 11928
rect 11978 11872 11980 11892
rect 11980 11872 12032 11892
rect 12032 11872 12034 11892
rect 11702 11348 11758 11384
rect 11702 11328 11704 11348
rect 11704 11328 11756 11348
rect 11756 11328 11758 11348
rect 11518 10784 11574 10840
rect 11518 10512 11574 10568
rect 11426 8628 11482 8664
rect 11426 8608 11428 8628
rect 11428 8608 11480 8628
rect 11480 8608 11482 8628
rect 11334 7384 11390 7440
rect 11334 7148 11336 7168
rect 11336 7148 11388 7168
rect 11388 7148 11390 7168
rect 11334 7112 11390 7148
rect 11610 8608 11666 8664
rect 11610 8084 11666 8120
rect 11610 8064 11612 8084
rect 11612 8064 11664 8084
rect 11664 8064 11666 8084
rect 11518 7520 11574 7576
rect 11426 6704 11482 6760
rect 10966 3984 11022 4040
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 12438 10920 12494 10976
rect 12438 10784 12494 10840
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 12438 10104 12494 10160
rect 12346 9832 12402 9888
rect 12254 9424 12310 9480
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 11978 8744 12034 8800
rect 12254 8900 12310 8936
rect 12254 8880 12256 8900
rect 12256 8880 12308 8900
rect 12308 8880 12310 8900
rect 12346 8744 12402 8800
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 11794 7656 11850 7712
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12714 13504 12770 13560
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 12806 12180 12808 12200
rect 12808 12180 12860 12200
rect 12860 12180 12862 12200
rect 12806 12144 12862 12180
rect 13082 15544 13138 15600
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12990 10512 13046 10568
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 13082 8472 13138 8528
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 11702 6432 11758 6488
rect 12622 7112 12678 7168
rect 12438 6568 12494 6624
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12714 6296 12770 6352
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 12530 5752 12586 5808
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 11702 3712 11758 3768
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12898 5888 12954 5944
rect 12898 5752 12954 5808
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12990 4140 13046 4176
rect 12990 4120 12992 4140
rect 12992 4120 13044 4140
rect 13044 4120 13046 4140
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 13726 17040 13782 17096
rect 14186 16652 14242 16688
rect 14186 16632 14188 16652
rect 14188 16632 14240 16652
rect 14240 16632 14242 16652
rect 13450 12280 13506 12336
rect 13910 13368 13966 13424
rect 13634 13252 13690 13288
rect 13634 13232 13636 13252
rect 13636 13232 13688 13252
rect 13688 13232 13690 13252
rect 13634 12008 13690 12064
rect 14094 13096 14150 13152
rect 13910 12708 13966 12744
rect 13910 12688 13912 12708
rect 13912 12688 13964 12708
rect 13964 12688 13966 12708
rect 13910 12552 13966 12608
rect 13818 11076 13874 11112
rect 13818 11056 13820 11076
rect 13820 11056 13872 11076
rect 13872 11056 13874 11076
rect 14094 11892 14150 11928
rect 14094 11872 14096 11892
rect 14096 11872 14148 11892
rect 14148 11872 14150 11892
rect 14094 11736 14150 11792
rect 13726 7792 13782 7848
rect 13634 7520 13690 7576
rect 14370 12180 14372 12200
rect 14372 12180 14424 12200
rect 14424 12180 14426 12200
rect 14370 12144 14426 12180
rect 14370 11872 14426 11928
rect 15290 13776 15346 13832
rect 14922 13096 14978 13152
rect 14922 12824 14978 12880
rect 13818 4800 13874 4856
rect 14370 8336 14426 8392
rect 15106 11736 15162 11792
rect 14278 6976 14334 7032
rect 14554 6860 14610 6896
rect 14554 6840 14556 6860
rect 14556 6840 14608 6860
rect 14608 6840 14610 6860
rect 14186 6296 14242 6352
rect 15198 11228 15200 11248
rect 15200 11228 15252 11248
rect 15252 11228 15254 11248
rect 15198 11192 15254 11228
rect 15198 9560 15254 9616
rect 14922 4548 14978 4584
rect 14922 4528 14924 4548
rect 14924 4528 14976 4548
rect 14976 4528 14978 4548
rect 15750 13812 15752 13832
rect 15752 13812 15804 13832
rect 15804 13812 15806 13832
rect 15750 13776 15806 13812
rect 15934 13912 15990 13968
rect 16118 13776 16174 13832
rect 15658 12280 15714 12336
rect 15658 11328 15714 11384
rect 15566 10648 15622 10704
rect 15382 7520 15438 7576
rect 15290 7112 15346 7168
rect 14922 2524 14924 2544
rect 14924 2524 14976 2544
rect 14976 2524 14978 2544
rect 14922 2488 14978 2524
rect 16026 11872 16082 11928
rect 16210 12552 16266 12608
rect 16118 6568 16174 6624
rect 16118 5208 16174 5264
rect 16026 4936 16082 4992
rect 16670 15408 16726 15464
rect 16670 12824 16726 12880
rect 16394 7384 16450 7440
rect 16578 12180 16580 12200
rect 16580 12180 16632 12200
rect 16632 12180 16634 12200
rect 16578 12144 16634 12180
rect 16578 11192 16634 11248
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 18510 16396 18512 16416
rect 18512 16396 18564 16416
rect 18564 16396 18566 16416
rect 18510 16360 18566 16396
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 17314 14320 17370 14376
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 18510 15308 18512 15328
rect 18512 15308 18564 15328
rect 18564 15308 18566 15328
rect 18510 15272 18566 15308
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 18234 14220 18236 14240
rect 18236 14220 18288 14240
rect 18288 14220 18290 14240
rect 18234 14184 18290 14220
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17038 11872 17094 11928
rect 17314 12044 17316 12064
rect 17316 12044 17368 12064
rect 17368 12044 17370 12064
rect 17314 12008 17370 12044
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16946 11192 17002 11248
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 17406 10920 17462 10976
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16854 6180 16910 6216
rect 16854 6160 16856 6180
rect 16856 6160 16908 6180
rect 16908 6160 16910 6180
rect 17314 6452 17370 6488
rect 17314 6432 17316 6452
rect 17316 6432 17368 6452
rect 17368 6432 17370 6452
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16854 5072 16910 5128
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 18510 13132 18512 13152
rect 18512 13132 18564 13152
rect 18564 13132 18566 13152
rect 18510 13096 18566 13132
rect 18050 6704 18106 6760
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 18510 12044 18512 12064
rect 18512 12044 18564 12064
rect 18564 12044 18566 12064
rect 18510 12008 18566 12044
rect 18326 11600 18382 11656
rect 18234 6316 18290 6352
rect 18234 6296 18236 6316
rect 18236 6296 18288 6316
rect 18288 6296 18290 6316
rect 18510 10920 18566 10976
rect 18510 9832 18566 9888
rect 18418 8880 18474 8936
rect 18418 8780 18420 8800
rect 18420 8780 18472 8800
rect 18472 8780 18474 8800
rect 18418 8744 18474 8780
rect 18418 7692 18420 7712
rect 18420 7692 18472 7712
rect 18472 7692 18474 7712
rect 18418 7656 18474 7692
rect 18418 6604 18420 6624
rect 18420 6604 18472 6624
rect 18472 6604 18474 6624
rect 18418 6568 18474 6604
rect 18418 5516 18420 5536
rect 18420 5516 18472 5536
rect 18472 5516 18474 5536
rect 18418 5480 18474 5516
rect 18234 4664 18290 4720
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 18418 4428 18420 4448
rect 18420 4428 18472 4448
rect 18472 4428 18474 4448
rect 18418 4392 18474 4428
rect 17866 3576 17922 3632
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 18418 3340 18420 3360
rect 18420 3340 18472 3360
rect 18472 3340 18474 3360
rect 18418 3304 18474 3340
rect 18142 3032 18198 3088
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 18786 12688 18842 12744
rect 18878 5616 18934 5672
rect 18418 2252 18420 2272
rect 18420 2252 18472 2272
rect 18472 2252 18474 2272
rect 18418 2216 18474 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
<< metal3 >>
rect 18505 17506 18571 17509
rect 19200 17506 20000 17536
rect 18505 17504 20000 17506
rect 18505 17448 18510 17504
rect 18566 17448 20000 17504
rect 18505 17446 20000 17448
rect 18505 17443 18571 17446
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 19200 17416 20000 17446
rect 17606 17375 17922 17376
rect 11605 17100 11671 17101
rect 11605 17098 11652 17100
rect 11564 17096 11652 17098
rect 11716 17098 11722 17100
rect 13721 17098 13787 17101
rect 11716 17096 13787 17098
rect 11564 17040 11610 17096
rect 11716 17040 13726 17096
rect 13782 17040 13787 17096
rect 11564 17038 11652 17040
rect 11605 17036 11652 17038
rect 11716 17038 13787 17040
rect 11716 17036 11722 17038
rect 11605 17035 11671 17036
rect 13721 17035 13787 17038
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 3325 16690 3391 16693
rect 14181 16690 14247 16693
rect 3325 16688 14247 16690
rect 3325 16632 3330 16688
rect 3386 16632 14186 16688
rect 14242 16632 14247 16688
rect 3325 16630 14247 16632
rect 3325 16627 3391 16630
rect 14181 16627 14247 16630
rect 18505 16418 18571 16421
rect 19200 16418 20000 16448
rect 18505 16416 20000 16418
rect 18505 16360 18510 16416
rect 18566 16360 20000 16416
rect 18505 16358 20000 16360
rect 18505 16355 18571 16358
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 19200 16328 20000 16358
rect 17606 16287 17922 16288
rect 8477 16010 8543 16013
rect 9438 16010 9444 16012
rect 8477 16008 9444 16010
rect 8477 15952 8482 16008
rect 8538 15952 9444 16008
rect 8477 15950 9444 15952
rect 8477 15947 8543 15950
rect 9438 15948 9444 15950
rect 9508 15948 9514 16012
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 5441 15602 5507 15605
rect 6361 15602 6427 15605
rect 5441 15600 6427 15602
rect 5441 15544 5446 15600
rect 5502 15544 6366 15600
rect 6422 15544 6427 15600
rect 5441 15542 6427 15544
rect 5441 15539 5507 15542
rect 6361 15539 6427 15542
rect 10317 15602 10383 15605
rect 13077 15602 13143 15605
rect 10317 15600 13143 15602
rect 10317 15544 10322 15600
rect 10378 15544 13082 15600
rect 13138 15544 13143 15600
rect 10317 15542 13143 15544
rect 10317 15539 10383 15542
rect 13077 15539 13143 15542
rect 4889 15466 4955 15469
rect 7833 15466 7899 15469
rect 16665 15466 16731 15469
rect 4889 15464 16731 15466
rect 4889 15408 4894 15464
rect 4950 15408 7838 15464
rect 7894 15408 16670 15464
rect 16726 15408 16731 15464
rect 4889 15406 16731 15408
rect 4889 15403 4955 15406
rect 7833 15403 7899 15406
rect 16665 15403 16731 15406
rect 1710 15268 1716 15332
rect 1780 15330 1786 15332
rect 2129 15330 2195 15333
rect 6085 15330 6151 15333
rect 1780 15328 2195 15330
rect 1780 15272 2134 15328
rect 2190 15272 2195 15328
rect 1780 15270 2195 15272
rect 1780 15268 1786 15270
rect 2129 15267 2195 15270
rect 3190 15328 6151 15330
rect 3190 15272 6090 15328
rect 6146 15272 6151 15328
rect 3190 15270 6151 15272
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 3190 15197 3250 15270
rect 6085 15267 6151 15270
rect 18505 15330 18571 15333
rect 19200 15330 20000 15360
rect 18505 15328 20000 15330
rect 18505 15272 18510 15328
rect 18566 15272 20000 15328
rect 18505 15270 20000 15272
rect 18505 15267 18571 15270
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 19200 15240 20000 15270
rect 17606 15199 17922 15200
rect 3141 15192 3250 15197
rect 3141 15136 3146 15192
rect 3202 15136 3250 15192
rect 3141 15134 3250 15136
rect 3141 15131 3207 15134
rect 0 15058 800 15088
rect 1577 15058 1643 15061
rect 0 15056 1643 15058
rect 0 15000 1582 15056
rect 1638 15000 1643 15056
rect 0 14998 1643 15000
rect 0 14968 800 14998
rect 1577 14995 1643 14998
rect 9305 15058 9371 15061
rect 10593 15058 10659 15061
rect 10869 15060 10935 15061
rect 10869 15058 10916 15060
rect 9305 15056 10659 15058
rect 9305 15000 9310 15056
rect 9366 15000 10598 15056
rect 10654 15000 10659 15056
rect 9305 14998 10659 15000
rect 10824 15056 10916 15058
rect 10824 15000 10874 15056
rect 10824 14998 10916 15000
rect 9305 14995 9371 14998
rect 10593 14995 10659 14998
rect 10869 14996 10916 14998
rect 10980 14996 10986 15060
rect 10869 14995 10935 14996
rect 10409 14922 10475 14925
rect 13670 14922 13676 14924
rect 10409 14920 13676 14922
rect 10409 14864 10414 14920
rect 10470 14864 13676 14920
rect 10409 14862 13676 14864
rect 10409 14859 10475 14862
rect 13670 14860 13676 14862
rect 13740 14860 13746 14924
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 5574 14452 5580 14516
rect 5644 14514 5650 14516
rect 10593 14514 10659 14517
rect 12433 14516 12499 14517
rect 12382 14514 12388 14516
rect 5644 14512 10659 14514
rect 5644 14456 10598 14512
rect 10654 14456 10659 14512
rect 5644 14454 10659 14456
rect 12342 14454 12388 14514
rect 12452 14512 12499 14516
rect 12494 14456 12499 14512
rect 5644 14452 5650 14454
rect 10593 14451 10659 14454
rect 12382 14452 12388 14454
rect 12452 14452 12499 14456
rect 12433 14451 12499 14452
rect 8109 14378 8175 14381
rect 17309 14378 17375 14381
rect 8109 14376 17375 14378
rect 8109 14320 8114 14376
rect 8170 14320 17314 14376
rect 17370 14320 17375 14376
rect 8109 14318 17375 14320
rect 8109 14315 8175 14318
rect 17309 14315 17375 14318
rect 18229 14242 18295 14245
rect 19200 14242 20000 14272
rect 18229 14240 20000 14242
rect 18229 14184 18234 14240
rect 18290 14184 20000 14240
rect 18229 14182 20000 14184
rect 18229 14179 18295 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 19200 14152 20000 14182
rect 17606 14111 17922 14112
rect 11094 14044 11100 14108
rect 11164 14106 11170 14108
rect 12065 14106 12131 14109
rect 11164 14104 12131 14106
rect 11164 14048 12070 14104
rect 12126 14048 12131 14104
rect 11164 14046 12131 14048
rect 11164 14044 11170 14046
rect 12065 14043 12131 14046
rect 4061 13970 4127 13973
rect 7557 13970 7623 13973
rect 4061 13968 7623 13970
rect 4061 13912 4066 13968
rect 4122 13912 7562 13968
rect 7618 13912 7623 13968
rect 4061 13910 7623 13912
rect 4061 13907 4127 13910
rect 7557 13907 7623 13910
rect 9622 13908 9628 13972
rect 9692 13970 9698 13972
rect 15929 13970 15995 13973
rect 9692 13968 15995 13970
rect 9692 13912 15934 13968
rect 15990 13912 15995 13968
rect 9692 13910 15995 13912
rect 9692 13908 9698 13910
rect 15929 13907 15995 13910
rect 6729 13836 6795 13837
rect 6678 13834 6684 13836
rect 6638 13774 6684 13834
rect 6748 13832 6795 13836
rect 6790 13776 6795 13832
rect 6678 13772 6684 13774
rect 6748 13772 6795 13776
rect 6729 13771 6795 13772
rect 10593 13834 10659 13837
rect 15285 13834 15351 13837
rect 10593 13832 15351 13834
rect 10593 13776 10598 13832
rect 10654 13776 15290 13832
rect 15346 13776 15351 13832
rect 10593 13774 15351 13776
rect 10593 13771 10659 13774
rect 15285 13771 15351 13774
rect 15510 13772 15516 13836
rect 15580 13834 15586 13836
rect 15745 13834 15811 13837
rect 15580 13832 15811 13834
rect 15580 13776 15750 13832
rect 15806 13776 15811 13832
rect 15580 13774 15811 13776
rect 15580 13772 15586 13774
rect 15745 13771 15811 13774
rect 16113 13834 16179 13837
rect 16246 13834 16252 13836
rect 16113 13832 16252 13834
rect 16113 13776 16118 13832
rect 16174 13776 16252 13832
rect 16113 13774 16252 13776
rect 16113 13771 16179 13774
rect 16246 13772 16252 13774
rect 16316 13772 16322 13836
rect 11462 13636 11468 13700
rect 11532 13698 11538 13700
rect 11789 13698 11855 13701
rect 11532 13696 11855 13698
rect 11532 13640 11794 13696
rect 11850 13640 11855 13696
rect 11532 13638 11855 13640
rect 11532 13636 11538 13638
rect 11789 13635 11855 13638
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 5625 13562 5691 13565
rect 2454 13560 5691 13562
rect 2454 13504 5630 13560
rect 5686 13504 5691 13560
rect 2454 13502 5691 13504
rect 1393 13426 1459 13429
rect 2454 13426 2514 13502
rect 5625 13499 5691 13502
rect 12709 13562 12775 13565
rect 13118 13562 13124 13564
rect 12709 13560 13124 13562
rect 12709 13504 12714 13560
rect 12770 13504 13124 13560
rect 12709 13502 13124 13504
rect 12709 13499 12775 13502
rect 13118 13500 13124 13502
rect 13188 13500 13194 13564
rect 1393 13424 2514 13426
rect 1393 13368 1398 13424
rect 1454 13368 2514 13424
rect 1393 13366 2514 13368
rect 4429 13426 4495 13429
rect 13905 13426 13971 13429
rect 4429 13424 13971 13426
rect 4429 13368 4434 13424
rect 4490 13368 13910 13424
rect 13966 13368 13971 13424
rect 4429 13366 13971 13368
rect 1393 13363 1459 13366
rect 4429 13363 4495 13366
rect 13905 13363 13971 13366
rect 2589 13290 2655 13293
rect 9949 13290 10015 13293
rect 10726 13290 10732 13292
rect 2589 13288 10732 13290
rect 2589 13232 2594 13288
rect 2650 13232 9954 13288
rect 10010 13232 10732 13288
rect 2589 13230 10732 13232
rect 2589 13227 2655 13230
rect 9949 13227 10015 13230
rect 10726 13228 10732 13230
rect 10796 13228 10802 13292
rect 13629 13290 13695 13293
rect 10872 13288 13695 13290
rect 10872 13232 13634 13288
rect 13690 13232 13695 13288
rect 10872 13230 13695 13232
rect 6545 13156 6611 13157
rect 6494 13154 6500 13156
rect 6454 13094 6500 13154
rect 6564 13152 6611 13156
rect 6606 13096 6611 13152
rect 6494 13092 6500 13094
rect 6564 13092 6611 13096
rect 6545 13091 6611 13092
rect 10225 13154 10291 13157
rect 10872 13154 10932 13230
rect 13629 13227 13695 13230
rect 10225 13152 10932 13154
rect 10225 13096 10230 13152
rect 10286 13096 10932 13152
rect 10225 13094 10932 13096
rect 14089 13154 14155 13157
rect 14222 13154 14228 13156
rect 14089 13152 14228 13154
rect 14089 13096 14094 13152
rect 14150 13096 14228 13152
rect 14089 13094 14228 13096
rect 10225 13091 10291 13094
rect 14089 13091 14155 13094
rect 14222 13092 14228 13094
rect 14292 13092 14298 13156
rect 14917 13154 14983 13157
rect 18505 13154 18571 13157
rect 19200 13154 20000 13184
rect 14917 13152 15026 13154
rect 14917 13096 14922 13152
rect 14978 13096 15026 13152
rect 14917 13091 15026 13096
rect 18505 13152 20000 13154
rect 18505 13096 18510 13152
rect 18566 13096 20000 13152
rect 18505 13094 20000 13096
rect 18505 13091 18571 13094
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 3693 13018 3759 13021
rect 7414 13018 7420 13020
rect 3693 13016 7420 13018
rect 3693 12960 3698 13016
rect 3754 12960 7420 13016
rect 3693 12958 7420 12960
rect 3693 12955 3759 12958
rect 7414 12956 7420 12958
rect 7484 12956 7490 13020
rect 10041 13018 10107 13021
rect 11145 13018 11211 13021
rect 10041 13016 11211 13018
rect 10041 12960 10046 13016
rect 10102 12960 11150 13016
rect 11206 12960 11211 13016
rect 10041 12958 11211 12960
rect 10041 12955 10107 12958
rect 11145 12955 11211 12958
rect 14966 12885 15026 13091
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 19200 13064 20000 13094
rect 17606 13023 17922 13024
rect 3918 12820 3924 12884
rect 3988 12882 3994 12884
rect 10961 12882 11027 12885
rect 3988 12880 11027 12882
rect 3988 12824 10966 12880
rect 11022 12824 11027 12880
rect 3988 12822 11027 12824
rect 3988 12820 3994 12822
rect 10961 12819 11027 12822
rect 14917 12880 15026 12885
rect 14917 12824 14922 12880
rect 14978 12824 15026 12880
rect 14917 12822 15026 12824
rect 16665 12882 16731 12885
rect 17350 12882 17356 12884
rect 16665 12880 17356 12882
rect 16665 12824 16670 12880
rect 16726 12824 17356 12880
rect 16665 12822 17356 12824
rect 14917 12819 14983 12822
rect 16665 12819 16731 12822
rect 17350 12820 17356 12822
rect 17420 12820 17426 12884
rect 1577 12746 1643 12749
rect 3049 12746 3115 12749
rect 13905 12746 13971 12749
rect 18781 12746 18847 12749
rect 1577 12744 2514 12746
rect 1577 12688 1582 12744
rect 1638 12688 2514 12744
rect 1577 12686 2514 12688
rect 1577 12683 1643 12686
rect 2454 12610 2514 12686
rect 3049 12744 12450 12746
rect 3049 12688 3054 12744
rect 3110 12688 12450 12744
rect 3049 12686 12450 12688
rect 3049 12683 3115 12686
rect 2454 12550 6746 12610
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6686 12338 6746 12550
rect 7414 12548 7420 12612
rect 7484 12610 7490 12612
rect 12390 12610 12450 12686
rect 13905 12744 18847 12746
rect 13905 12688 13910 12744
rect 13966 12688 18786 12744
rect 18842 12688 18847 12744
rect 13905 12686 18847 12688
rect 13905 12683 13971 12686
rect 18781 12683 18847 12686
rect 13905 12610 13971 12613
rect 7484 12550 11714 12610
rect 12390 12608 13971 12610
rect 12390 12552 13910 12608
rect 13966 12552 13971 12608
rect 12390 12550 13971 12552
rect 7484 12548 7490 12550
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 8569 12474 8635 12477
rect 7422 12472 8635 12474
rect 7422 12416 8574 12472
rect 8630 12416 8635 12472
rect 7422 12414 8635 12416
rect 7422 12338 7482 12414
rect 8569 12411 8635 12414
rect 6686 12278 7482 12338
rect 11654 12338 11714 12550
rect 13905 12547 13971 12550
rect 15142 12548 15148 12612
rect 15212 12610 15218 12612
rect 16205 12610 16271 12613
rect 15212 12608 16271 12610
rect 15212 12552 16210 12608
rect 16266 12552 16271 12608
rect 15212 12550 16271 12552
rect 15212 12548 15218 12550
rect 16205 12547 16271 12550
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 13302 12338 13308 12340
rect 11654 12278 13308 12338
rect 13302 12276 13308 12278
rect 13372 12276 13378 12340
rect 13445 12338 13511 12341
rect 15653 12338 15719 12341
rect 13445 12336 15719 12338
rect 13445 12280 13450 12336
rect 13506 12280 15658 12336
rect 15714 12280 15719 12336
rect 13445 12278 15719 12280
rect 13445 12275 13511 12278
rect 15653 12275 15719 12278
rect 4705 12202 4771 12205
rect 8293 12202 8359 12205
rect 12801 12202 12867 12205
rect 4705 12200 12867 12202
rect 4705 12144 4710 12200
rect 4766 12144 8298 12200
rect 8354 12144 12806 12200
rect 12862 12144 12867 12200
rect 4705 12142 12867 12144
rect 4705 12139 4771 12142
rect 8293 12139 8359 12142
rect 12801 12139 12867 12142
rect 14365 12202 14431 12205
rect 16573 12202 16639 12205
rect 14365 12200 16639 12202
rect 14365 12144 14370 12200
rect 14426 12144 16578 12200
rect 16634 12144 16639 12200
rect 14365 12142 16639 12144
rect 14365 12139 14431 12142
rect 16573 12139 16639 12142
rect 6821 12066 6887 12069
rect 7414 12066 7420 12068
rect 6821 12064 7420 12066
rect 6821 12008 6826 12064
rect 6882 12008 7420 12064
rect 6821 12006 7420 12008
rect 6821 12003 6887 12006
rect 7414 12004 7420 12006
rect 7484 12004 7490 12068
rect 13629 12066 13695 12069
rect 17309 12066 17375 12069
rect 13629 12064 17375 12066
rect 13629 12008 13634 12064
rect 13690 12008 17314 12064
rect 17370 12008 17375 12064
rect 13629 12006 17375 12008
rect 13629 12003 13695 12006
rect 17309 12003 17375 12006
rect 18505 12066 18571 12069
rect 19200 12066 20000 12096
rect 18505 12064 20000 12066
rect 18505 12008 18510 12064
rect 18566 12008 20000 12064
rect 18505 12006 20000 12008
rect 18505 12003 18571 12006
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 19200 11976 20000 12006
rect 17606 11935 17922 11936
rect 6545 11930 6611 11933
rect 7465 11930 7531 11933
rect 6545 11928 7531 11930
rect 6545 11872 6550 11928
rect 6606 11872 7470 11928
rect 7526 11872 7531 11928
rect 6545 11870 7531 11872
rect 6545 11867 6611 11870
rect 7465 11867 7531 11870
rect 8661 11930 8727 11933
rect 9489 11930 9555 11933
rect 9949 11932 10015 11933
rect 9949 11930 9996 11932
rect 8661 11928 9555 11930
rect 8661 11872 8666 11928
rect 8722 11872 9494 11928
rect 9550 11872 9555 11928
rect 8661 11870 9555 11872
rect 9904 11928 9996 11930
rect 9904 11872 9954 11928
rect 9904 11870 9996 11872
rect 8661 11867 8727 11870
rect 9489 11867 9555 11870
rect 9949 11868 9996 11870
rect 10060 11868 10066 11932
rect 10593 11930 10659 11933
rect 11973 11930 12039 11933
rect 10593 11928 12039 11930
rect 10593 11872 10598 11928
rect 10654 11872 11978 11928
rect 12034 11872 12039 11928
rect 10593 11870 12039 11872
rect 9949 11867 10015 11868
rect 10593 11867 10659 11870
rect 11973 11867 12039 11870
rect 13854 11868 13860 11932
rect 13924 11930 13930 11932
rect 14089 11930 14155 11933
rect 13924 11928 14155 11930
rect 13924 11872 14094 11928
rect 14150 11872 14155 11928
rect 13924 11870 14155 11872
rect 13924 11868 13930 11870
rect 14089 11867 14155 11870
rect 14365 11930 14431 11933
rect 16021 11930 16087 11933
rect 14365 11928 16087 11930
rect 14365 11872 14370 11928
rect 14426 11872 16026 11928
rect 16082 11872 16087 11928
rect 14365 11870 16087 11872
rect 14365 11867 14431 11870
rect 16021 11867 16087 11870
rect 16614 11868 16620 11932
rect 16684 11930 16690 11932
rect 17033 11930 17099 11933
rect 16684 11928 17099 11930
rect 16684 11872 17038 11928
rect 17094 11872 17099 11928
rect 16684 11870 17099 11872
rect 16684 11868 16690 11870
rect 17033 11867 17099 11870
rect 4521 11794 4587 11797
rect 7741 11794 7807 11797
rect 4521 11792 7807 11794
rect 4521 11736 4526 11792
rect 4582 11736 7746 11792
rect 7802 11736 7807 11792
rect 4521 11734 7807 11736
rect 4521 11731 4587 11734
rect 7741 11731 7807 11734
rect 7925 11794 7991 11797
rect 14089 11794 14155 11797
rect 15101 11794 15167 11797
rect 7925 11792 15167 11794
rect 7925 11736 7930 11792
rect 7986 11736 14094 11792
rect 14150 11736 15106 11792
rect 15162 11736 15167 11792
rect 7925 11734 15167 11736
rect 7925 11731 7991 11734
rect 14089 11731 14155 11734
rect 15101 11731 15167 11734
rect 5625 11658 5691 11661
rect 18321 11658 18387 11661
rect 5625 11656 18387 11658
rect 5625 11600 5630 11656
rect 5686 11600 18326 11656
rect 18382 11600 18387 11656
rect 5625 11598 18387 11600
rect 5625 11595 5691 11598
rect 18321 11595 18387 11598
rect 3693 11524 3759 11525
rect 3693 11522 3740 11524
rect 3648 11520 3740 11522
rect 3648 11464 3698 11520
rect 3648 11462 3740 11464
rect 3693 11460 3740 11462
rect 3804 11460 3810 11524
rect 7741 11522 7807 11525
rect 8518 11522 8524 11524
rect 7741 11520 8524 11522
rect 7741 11464 7746 11520
rect 7802 11464 8524 11520
rect 7741 11462 8524 11464
rect 3693 11459 3759 11460
rect 7741 11459 7807 11462
rect 8518 11460 8524 11462
rect 8588 11460 8594 11524
rect 10910 11460 10916 11524
rect 10980 11522 10986 11524
rect 11329 11522 11395 11525
rect 10980 11520 11395 11522
rect 10980 11464 11334 11520
rect 11390 11464 11395 11520
rect 10980 11462 11395 11464
rect 10980 11460 10986 11462
rect 11329 11459 11395 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 9990 11324 9996 11388
rect 10060 11386 10066 11388
rect 11145 11386 11211 11389
rect 11697 11388 11763 11389
rect 10060 11384 11211 11386
rect 10060 11328 11150 11384
rect 11206 11328 11211 11384
rect 10060 11326 11211 11328
rect 10060 11324 10066 11326
rect 11145 11323 11211 11326
rect 11646 11324 11652 11388
rect 11716 11386 11763 11388
rect 11716 11384 11808 11386
rect 11758 11328 11808 11384
rect 11716 11326 11808 11328
rect 11716 11324 11763 11326
rect 14038 11324 14044 11388
rect 14108 11386 14114 11388
rect 15653 11386 15719 11389
rect 14108 11384 15719 11386
rect 14108 11328 15658 11384
rect 15714 11328 15719 11384
rect 14108 11326 15719 11328
rect 14108 11324 14114 11326
rect 11697 11323 11763 11324
rect 15653 11323 15719 11326
rect 7741 11250 7807 11253
rect 9305 11250 9371 11253
rect 7741 11248 9371 11250
rect 7741 11192 7746 11248
rect 7802 11192 9310 11248
rect 9366 11192 9371 11248
rect 7741 11190 9371 11192
rect 7741 11187 7807 11190
rect 9305 11187 9371 11190
rect 9673 11250 9739 11253
rect 15193 11250 15259 11253
rect 9673 11248 15259 11250
rect 9673 11192 9678 11248
rect 9734 11192 15198 11248
rect 15254 11192 15259 11248
rect 9673 11190 15259 11192
rect 9673 11187 9739 11190
rect 15193 11187 15259 11190
rect 16573 11250 16639 11253
rect 16941 11250 17007 11253
rect 16573 11248 17007 11250
rect 16573 11192 16578 11248
rect 16634 11192 16946 11248
rect 17002 11192 17007 11248
rect 16573 11190 17007 11192
rect 16573 11187 16639 11190
rect 16941 11187 17007 11190
rect 10501 11114 10567 11117
rect 11646 11114 11652 11116
rect 10501 11112 11652 11114
rect 10501 11056 10506 11112
rect 10562 11056 11652 11112
rect 10501 11054 11652 11056
rect 10501 11051 10567 11054
rect 11646 11052 11652 11054
rect 11716 11052 11722 11116
rect 13670 11052 13676 11116
rect 13740 11114 13746 11116
rect 13813 11114 13879 11117
rect 13740 11112 13879 11114
rect 13740 11056 13818 11112
rect 13874 11056 13879 11112
rect 13740 11054 13879 11056
rect 13740 11052 13746 11054
rect 13813 11051 13879 11054
rect 9397 10978 9463 10981
rect 9622 10978 9628 10980
rect 9397 10976 9628 10978
rect 9397 10920 9402 10976
rect 9458 10920 9628 10976
rect 9397 10918 9628 10920
rect 9397 10915 9463 10918
rect 9622 10916 9628 10918
rect 9692 10916 9698 10980
rect 11237 10978 11303 10981
rect 12433 10978 12499 10981
rect 17401 10980 17467 10981
rect 11237 10976 12499 10978
rect 11237 10920 11242 10976
rect 11298 10920 12438 10976
rect 12494 10920 12499 10976
rect 11237 10918 12499 10920
rect 11237 10915 11303 10918
rect 12433 10915 12499 10918
rect 17350 10916 17356 10980
rect 17420 10978 17467 10980
rect 18505 10978 18571 10981
rect 19200 10978 20000 11008
rect 17420 10976 17512 10978
rect 17462 10920 17512 10976
rect 17420 10918 17512 10920
rect 18505 10976 20000 10978
rect 18505 10920 18510 10976
rect 18566 10920 20000 10976
rect 18505 10918 20000 10920
rect 17420 10916 17467 10918
rect 17401 10915 17467 10916
rect 18505 10915 18571 10918
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 19200 10888 20000 10918
rect 17606 10847 17922 10848
rect 9581 10844 9647 10845
rect 9581 10840 9628 10844
rect 9692 10842 9698 10844
rect 9581 10784 9586 10840
rect 9581 10780 9628 10784
rect 9692 10782 9738 10842
rect 9692 10780 9698 10782
rect 11094 10780 11100 10844
rect 11164 10842 11170 10844
rect 11329 10842 11395 10845
rect 11164 10840 11395 10842
rect 11164 10784 11334 10840
rect 11390 10784 11395 10840
rect 11164 10782 11395 10784
rect 11164 10780 11170 10782
rect 9581 10779 9647 10780
rect 11329 10779 11395 10782
rect 11513 10842 11579 10845
rect 12433 10844 12499 10845
rect 11646 10842 11652 10844
rect 11513 10840 11652 10842
rect 11513 10784 11518 10840
rect 11574 10784 11652 10840
rect 11513 10782 11652 10784
rect 11513 10779 11579 10782
rect 11646 10780 11652 10782
rect 11716 10780 11722 10844
rect 12382 10780 12388 10844
rect 12452 10842 12499 10844
rect 12452 10840 12544 10842
rect 12494 10784 12544 10840
rect 12452 10782 12544 10784
rect 12452 10780 12499 10782
rect 12433 10779 12499 10780
rect 2589 10706 2655 10709
rect 15561 10706 15627 10709
rect 2589 10704 15627 10706
rect 2589 10648 2594 10704
rect 2650 10648 15566 10704
rect 15622 10648 15627 10704
rect 2589 10646 15627 10648
rect 2589 10643 2655 10646
rect 15561 10643 15627 10646
rect 4061 10570 4127 10573
rect 8334 10570 8340 10572
rect 4061 10568 8340 10570
rect 4061 10512 4066 10568
rect 4122 10512 8340 10568
rect 4061 10510 8340 10512
rect 4061 10507 4127 10510
rect 8334 10508 8340 10510
rect 8404 10508 8410 10572
rect 11513 10570 11579 10573
rect 12985 10570 13051 10573
rect 11513 10568 13051 10570
rect 11513 10512 11518 10568
rect 11574 10512 12990 10568
rect 13046 10512 13051 10568
rect 11513 10510 13051 10512
rect 11513 10507 11579 10510
rect 12985 10507 13051 10510
rect 8569 10434 8635 10437
rect 8702 10434 8708 10436
rect 8569 10432 8708 10434
rect 8569 10376 8574 10432
rect 8630 10376 8708 10432
rect 8569 10374 8708 10376
rect 8569 10371 8635 10374
rect 8702 10372 8708 10374
rect 8772 10372 8778 10436
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 8661 10298 8727 10301
rect 8886 10298 8892 10300
rect 8661 10296 8892 10298
rect 8661 10240 8666 10296
rect 8722 10240 8892 10296
rect 8661 10238 8892 10240
rect 8661 10235 8727 10238
rect 8886 10236 8892 10238
rect 8956 10236 8962 10300
rect 4337 10162 4403 10165
rect 12433 10162 12499 10165
rect 4337 10160 12499 10162
rect 4337 10104 4342 10160
rect 4398 10104 12438 10160
rect 12494 10104 12499 10160
rect 4337 10102 12499 10104
rect 4337 10099 4403 10102
rect 12433 10099 12499 10102
rect 5390 9964 5396 10028
rect 5460 10026 5466 10028
rect 8661 10026 8727 10029
rect 5460 10024 8727 10026
rect 5460 9968 8666 10024
rect 8722 9968 8727 10024
rect 5460 9966 8727 9968
rect 5460 9964 5466 9966
rect 8661 9963 8727 9966
rect 9581 9890 9647 9893
rect 12341 9890 12407 9893
rect 9581 9888 12407 9890
rect 9581 9832 9586 9888
rect 9642 9832 12346 9888
rect 12402 9832 12407 9888
rect 9581 9830 12407 9832
rect 9581 9827 9647 9830
rect 12341 9827 12407 9830
rect 18505 9890 18571 9893
rect 19200 9890 20000 9920
rect 18505 9888 20000 9890
rect 18505 9832 18510 9888
rect 18566 9832 20000 9888
rect 18505 9830 20000 9832
rect 18505 9827 18571 9830
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 19200 9800 20000 9830
rect 17606 9759 17922 9760
rect 3049 9754 3115 9757
rect 5574 9754 5580 9756
rect 3049 9752 5580 9754
rect 3049 9696 3054 9752
rect 3110 9696 5580 9752
rect 3049 9694 5580 9696
rect 3049 9691 3115 9694
rect 5574 9692 5580 9694
rect 5644 9692 5650 9756
rect 6361 9754 6427 9757
rect 6678 9754 6684 9756
rect 6361 9752 6684 9754
rect 6361 9696 6366 9752
rect 6422 9696 6684 9752
rect 6361 9694 6684 9696
rect 6361 9691 6427 9694
rect 6678 9692 6684 9694
rect 6748 9692 6754 9756
rect 8569 9754 8635 9757
rect 9489 9754 9555 9757
rect 10542 9754 10548 9756
rect 8569 9752 9555 9754
rect 8569 9696 8574 9752
rect 8630 9696 9494 9752
rect 9550 9696 9555 9752
rect 8569 9694 9555 9696
rect 8569 9691 8635 9694
rect 9489 9691 9555 9694
rect 10366 9694 10548 9754
rect 1669 9618 1735 9621
rect 4521 9618 4587 9621
rect 1669 9616 4587 9618
rect 1669 9560 1674 9616
rect 1730 9560 4526 9616
rect 4582 9560 4587 9616
rect 1669 9558 4587 9560
rect 1669 9555 1735 9558
rect 4521 9555 4587 9558
rect 5993 9618 6059 9621
rect 6821 9618 6887 9621
rect 10366 9618 10426 9694
rect 10542 9692 10548 9694
rect 10612 9754 10618 9756
rect 10961 9754 11027 9757
rect 10612 9752 11027 9754
rect 10612 9696 10966 9752
rect 11022 9696 11027 9752
rect 10612 9694 11027 9696
rect 10612 9692 10618 9694
rect 10961 9691 11027 9694
rect 5993 9616 10426 9618
rect 5993 9560 5998 9616
rect 6054 9560 6826 9616
rect 6882 9560 10426 9616
rect 5993 9558 10426 9560
rect 11237 9618 11303 9621
rect 15193 9618 15259 9621
rect 11237 9616 15259 9618
rect 11237 9560 11242 9616
rect 11298 9560 15198 9616
rect 15254 9560 15259 9616
rect 11237 9558 15259 9560
rect 5993 9555 6059 9558
rect 6821 9555 6887 9558
rect 11237 9555 11303 9558
rect 15193 9555 15259 9558
rect 2405 9482 2471 9485
rect 9806 9482 9812 9484
rect 2405 9480 9812 9482
rect 2405 9424 2410 9480
rect 2466 9424 9812 9480
rect 2405 9422 9812 9424
rect 2405 9419 2471 9422
rect 9806 9420 9812 9422
rect 9876 9420 9882 9484
rect 11278 9420 11284 9484
rect 11348 9482 11354 9484
rect 12249 9482 12315 9485
rect 11348 9480 12315 9482
rect 11348 9424 12254 9480
rect 12310 9424 12315 9480
rect 11348 9422 12315 9424
rect 11348 9420 11354 9422
rect 12249 9419 12315 9422
rect 7741 9346 7807 9349
rect 8150 9346 8156 9348
rect 7741 9344 8156 9346
rect 7741 9288 7746 9344
rect 7802 9288 8156 9344
rect 7741 9286 8156 9288
rect 7741 9283 7807 9286
rect 8150 9284 8156 9286
rect 8220 9284 8226 9348
rect 9070 9284 9076 9348
rect 9140 9346 9146 9348
rect 9397 9346 9463 9349
rect 9140 9344 9463 9346
rect 9140 9288 9402 9344
rect 9458 9288 9463 9344
rect 9140 9286 9463 9288
rect 9140 9284 9146 9286
rect 9397 9283 9463 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 7925 9210 7991 9213
rect 8886 9210 8892 9212
rect 7925 9208 8892 9210
rect 7925 9152 7930 9208
rect 7986 9152 8892 9208
rect 7925 9150 8892 9152
rect 7925 9147 7991 9150
rect 8886 9148 8892 9150
rect 8956 9210 8962 9212
rect 10685 9210 10751 9213
rect 8956 9208 10751 9210
rect 8956 9152 10690 9208
rect 10746 9152 10751 9208
rect 8956 9150 10751 9152
rect 8956 9148 8962 9150
rect 10685 9147 10751 9150
rect 4337 9074 4403 9077
rect 13854 9074 13860 9076
rect 4337 9072 13860 9074
rect 4337 9016 4342 9072
rect 4398 9016 13860 9072
rect 4337 9014 13860 9016
rect 4337 9011 4403 9014
rect 13854 9012 13860 9014
rect 13924 9012 13930 9076
rect 4061 8938 4127 8941
rect 6269 8938 6335 8941
rect 8150 8938 8156 8940
rect 4061 8936 8156 8938
rect 4061 8880 4066 8936
rect 4122 8880 6274 8936
rect 6330 8880 8156 8936
rect 4061 8878 8156 8880
rect 4061 8875 4127 8878
rect 6269 8875 6335 8878
rect 8150 8876 8156 8878
rect 8220 8938 8226 8940
rect 8569 8938 8635 8941
rect 8220 8936 8635 8938
rect 8220 8880 8574 8936
rect 8630 8880 8635 8936
rect 8220 8878 8635 8880
rect 8220 8876 8226 8878
rect 8569 8875 8635 8878
rect 9213 8938 9279 8941
rect 10409 8938 10475 8941
rect 9213 8936 10475 8938
rect 9213 8880 9218 8936
rect 9274 8880 10414 8936
rect 10470 8880 10475 8936
rect 9213 8878 10475 8880
rect 9213 8875 9279 8878
rect 10409 8875 10475 8878
rect 11145 8938 11211 8941
rect 12249 8938 12315 8941
rect 17350 8938 17356 8940
rect 11145 8936 12315 8938
rect 11145 8880 11150 8936
rect 11206 8880 12254 8936
rect 12310 8880 12315 8936
rect 11145 8878 12315 8880
rect 11145 8875 11211 8878
rect 12249 8875 12315 8878
rect 12390 8878 17356 8938
rect 12390 8805 12450 8878
rect 17350 8876 17356 8878
rect 17420 8938 17426 8940
rect 18413 8938 18479 8941
rect 17420 8936 18479 8938
rect 17420 8880 18418 8936
rect 18474 8880 18479 8936
rect 17420 8878 18479 8880
rect 17420 8876 17426 8878
rect 18413 8875 18479 8878
rect 5993 8802 6059 8805
rect 6269 8802 6335 8805
rect 5993 8800 6335 8802
rect 5993 8744 5998 8800
rect 6054 8744 6274 8800
rect 6330 8744 6335 8800
rect 5993 8742 6335 8744
rect 5993 8739 6059 8742
rect 6269 8739 6335 8742
rect 8334 8740 8340 8804
rect 8404 8802 8410 8804
rect 8477 8802 8543 8805
rect 8404 8800 8543 8802
rect 8404 8744 8482 8800
rect 8538 8744 8543 8800
rect 8404 8742 8543 8744
rect 8404 8740 8410 8742
rect 8477 8739 8543 8742
rect 10133 8802 10199 8805
rect 10409 8802 10475 8805
rect 10133 8800 10475 8802
rect 10133 8744 10138 8800
rect 10194 8744 10414 8800
rect 10470 8744 10475 8800
rect 10133 8742 10475 8744
rect 10133 8739 10199 8742
rect 10409 8739 10475 8742
rect 10685 8802 10751 8805
rect 11973 8802 12039 8805
rect 10685 8800 12039 8802
rect 10685 8744 10690 8800
rect 10746 8744 11978 8800
rect 12034 8744 12039 8800
rect 10685 8742 12039 8744
rect 10685 8739 10751 8742
rect 11973 8739 12039 8742
rect 12341 8800 12450 8805
rect 12341 8744 12346 8800
rect 12402 8744 12450 8800
rect 12341 8742 12450 8744
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 12341 8739 12407 8742
rect 18413 8739 18479 8742
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 19200 8712 20000 8742
rect 17606 8671 17922 8672
rect 4061 8666 4127 8669
rect 4245 8666 4311 8669
rect 4061 8664 4311 8666
rect 4061 8608 4066 8664
rect 4122 8608 4250 8664
rect 4306 8608 4311 8664
rect 4061 8606 4311 8608
rect 4061 8603 4127 8606
rect 4245 8603 4311 8606
rect 8661 8666 8727 8669
rect 11421 8666 11487 8669
rect 8661 8664 11487 8666
rect 8661 8608 8666 8664
rect 8722 8608 11426 8664
rect 11482 8608 11487 8664
rect 8661 8606 11487 8608
rect 8661 8603 8727 8606
rect 11421 8603 11487 8606
rect 11605 8666 11671 8669
rect 11605 8664 12496 8666
rect 11605 8608 11610 8664
rect 11666 8608 12496 8664
rect 11605 8606 12496 8608
rect 11605 8603 11671 8606
rect 4153 8530 4219 8533
rect 11237 8530 11303 8533
rect 4153 8528 11303 8530
rect 4153 8472 4158 8528
rect 4214 8472 11242 8528
rect 11298 8472 11303 8528
rect 4153 8470 11303 8472
rect 12436 8530 12496 8606
rect 13077 8530 13143 8533
rect 12436 8528 13143 8530
rect 12436 8472 13082 8528
rect 13138 8472 13143 8528
rect 12436 8470 13143 8472
rect 4153 8467 4219 8470
rect 11237 8467 11303 8470
rect 13077 8467 13143 8470
rect 1945 8394 2011 8397
rect 4245 8394 4311 8397
rect 4797 8394 4863 8397
rect 1945 8392 4863 8394
rect 1945 8336 1950 8392
rect 2006 8336 4250 8392
rect 4306 8336 4802 8392
rect 4858 8336 4863 8392
rect 1945 8334 4863 8336
rect 1945 8331 2011 8334
rect 4245 8331 4311 8334
rect 4797 8331 4863 8334
rect 5349 8394 5415 8397
rect 9121 8394 9187 8397
rect 5349 8392 9187 8394
rect 5349 8336 5354 8392
rect 5410 8336 9126 8392
rect 9182 8336 9187 8392
rect 5349 8334 9187 8336
rect 5349 8331 5415 8334
rect 9121 8331 9187 8334
rect 9673 8394 9739 8397
rect 11237 8394 11303 8397
rect 14365 8394 14431 8397
rect 9673 8392 11303 8394
rect 9673 8336 9678 8392
rect 9734 8336 11242 8392
rect 11298 8336 11303 8392
rect 9673 8334 11303 8336
rect 9673 8331 9739 8334
rect 11237 8331 11303 8334
rect 11654 8392 14431 8394
rect 11654 8336 14370 8392
rect 14426 8336 14431 8392
rect 11654 8334 14431 8336
rect 3509 8258 3575 8261
rect 5717 8258 5783 8261
rect 3509 8256 5783 8258
rect 3509 8200 3514 8256
rect 3570 8200 5722 8256
rect 5778 8200 5783 8256
rect 3509 8198 5783 8200
rect 3509 8195 3575 8198
rect 5717 8195 5783 8198
rect 8661 8260 8727 8261
rect 8661 8256 8708 8260
rect 8772 8258 8778 8260
rect 10225 8258 10291 8261
rect 11654 8258 11714 8334
rect 14365 8331 14431 8334
rect 8661 8200 8666 8256
rect 8661 8196 8708 8200
rect 8772 8198 8818 8258
rect 10225 8256 11714 8258
rect 10225 8200 10230 8256
rect 10286 8200 11714 8256
rect 10225 8198 11714 8200
rect 8772 8196 8778 8198
rect 8661 8195 8727 8196
rect 10225 8195 10291 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 7557 8122 7623 8125
rect 9070 8122 9076 8124
rect 7557 8120 9076 8122
rect 7557 8064 7562 8120
rect 7618 8064 9076 8120
rect 7557 8062 9076 8064
rect 7557 8059 7623 8062
rect 9070 8060 9076 8062
rect 9140 8060 9146 8124
rect 9673 8122 9739 8125
rect 11605 8122 11671 8125
rect 9673 8120 11671 8122
rect 9673 8064 9678 8120
rect 9734 8064 11610 8120
rect 11666 8064 11671 8120
rect 9673 8062 11671 8064
rect 9673 8059 9739 8062
rect 11605 8059 11671 8062
rect 3877 7986 3943 7989
rect 9489 7986 9555 7989
rect 3877 7984 9555 7986
rect 3877 7928 3882 7984
rect 3938 7928 9494 7984
rect 9550 7928 9555 7984
rect 3877 7926 9555 7928
rect 3877 7923 3943 7926
rect 9489 7923 9555 7926
rect 11053 7986 11119 7989
rect 14038 7986 14044 7988
rect 11053 7984 14044 7986
rect 11053 7928 11058 7984
rect 11114 7928 14044 7984
rect 11053 7926 14044 7928
rect 11053 7923 11119 7926
rect 14038 7924 14044 7926
rect 14108 7924 14114 7988
rect 3877 7850 3943 7853
rect 5901 7850 5967 7853
rect 3877 7848 5967 7850
rect 3877 7792 3882 7848
rect 3938 7792 5906 7848
rect 5962 7792 5967 7848
rect 3877 7790 5967 7792
rect 3877 7787 3943 7790
rect 5901 7787 5967 7790
rect 6085 7850 6151 7853
rect 7557 7850 7623 7853
rect 6085 7848 7623 7850
rect 6085 7792 6090 7848
rect 6146 7792 7562 7848
rect 7618 7792 7623 7848
rect 6085 7790 7623 7792
rect 6085 7787 6151 7790
rect 7557 7787 7623 7790
rect 7833 7850 7899 7853
rect 11053 7850 11119 7853
rect 7833 7848 11119 7850
rect 7833 7792 7838 7848
rect 7894 7792 11058 7848
rect 11114 7792 11119 7848
rect 7833 7790 11119 7792
rect 7833 7787 7899 7790
rect 11053 7787 11119 7790
rect 11462 7788 11468 7852
rect 11532 7850 11538 7852
rect 13721 7850 13787 7853
rect 11532 7848 13787 7850
rect 11532 7792 13726 7848
rect 13782 7792 13787 7848
rect 11532 7790 13787 7792
rect 11532 7788 11538 7790
rect 13721 7787 13787 7790
rect 11094 7652 11100 7716
rect 11164 7714 11170 7716
rect 11789 7714 11855 7717
rect 11164 7712 11855 7714
rect 11164 7656 11794 7712
rect 11850 7656 11855 7712
rect 11164 7654 11855 7656
rect 11164 7652 11170 7654
rect 11789 7651 11855 7654
rect 18413 7714 18479 7717
rect 19200 7714 20000 7744
rect 18413 7712 20000 7714
rect 18413 7656 18418 7712
rect 18474 7656 20000 7712
rect 18413 7654 20000 7656
rect 18413 7651 18479 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 19200 7624 20000 7654
rect 17606 7583 17922 7584
rect 10542 7516 10548 7580
rect 10612 7578 10618 7580
rect 11513 7578 11579 7581
rect 10612 7576 11579 7578
rect 10612 7520 11518 7576
rect 11574 7520 11579 7576
rect 10612 7518 11579 7520
rect 10612 7516 10618 7518
rect 11513 7515 11579 7518
rect 13629 7578 13695 7581
rect 15377 7578 15443 7581
rect 13629 7576 15443 7578
rect 13629 7520 13634 7576
rect 13690 7520 15382 7576
rect 15438 7520 15443 7576
rect 13629 7518 15443 7520
rect 13629 7515 13695 7518
rect 15377 7515 15443 7518
rect 2681 7442 2747 7445
rect 3049 7442 3115 7445
rect 2681 7440 3115 7442
rect 2681 7384 2686 7440
rect 2742 7384 3054 7440
rect 3110 7384 3115 7440
rect 2681 7382 3115 7384
rect 2681 7379 2747 7382
rect 3049 7379 3115 7382
rect 6361 7442 6427 7445
rect 11329 7442 11395 7445
rect 16389 7442 16455 7445
rect 6361 7440 16455 7442
rect 6361 7384 6366 7440
rect 6422 7384 11334 7440
rect 11390 7384 16394 7440
rect 16450 7384 16455 7440
rect 6361 7382 16455 7384
rect 6361 7379 6427 7382
rect 11329 7379 11395 7382
rect 16389 7379 16455 7382
rect 5901 7306 5967 7309
rect 15142 7306 15148 7308
rect 5901 7304 15148 7306
rect 5901 7248 5906 7304
rect 5962 7248 15148 7304
rect 5901 7246 15148 7248
rect 5901 7243 5967 7246
rect 15142 7244 15148 7246
rect 15212 7244 15218 7308
rect 11329 7172 11395 7173
rect 11278 7108 11284 7172
rect 11348 7170 11395 7172
rect 12617 7170 12683 7173
rect 15285 7170 15351 7173
rect 11348 7168 11440 7170
rect 11390 7112 11440 7168
rect 11348 7110 11440 7112
rect 12617 7168 15351 7170
rect 12617 7112 12622 7168
rect 12678 7112 15290 7168
rect 15346 7112 15351 7168
rect 12617 7110 15351 7112
rect 11348 7108 11395 7110
rect 11329 7107 11395 7108
rect 12617 7107 12683 7110
rect 15285 7107 15351 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 3509 7034 3575 7037
rect 11462 7034 11468 7036
rect 3509 7032 6746 7034
rect 3509 6976 3514 7032
rect 3570 6976 6746 7032
rect 3509 6974 6746 6976
rect 3509 6971 3575 6974
rect 6686 6898 6746 6974
rect 7422 6974 11468 7034
rect 7422 6898 7482 6974
rect 11462 6972 11468 6974
rect 11532 6972 11538 7036
rect 13302 6972 13308 7036
rect 13372 7034 13378 7036
rect 14273 7034 14339 7037
rect 13372 7032 14339 7034
rect 13372 6976 14278 7032
rect 14334 6976 14339 7032
rect 13372 6974 14339 6976
rect 13372 6972 13378 6974
rect 14273 6971 14339 6974
rect 6686 6838 7482 6898
rect 9806 6836 9812 6900
rect 9876 6898 9882 6900
rect 14549 6898 14615 6901
rect 9876 6896 14615 6898
rect 9876 6840 14554 6896
rect 14610 6840 14615 6896
rect 9876 6838 14615 6840
rect 9876 6836 9882 6838
rect 14549 6835 14615 6838
rect 4797 6764 4863 6765
rect 4797 6762 4844 6764
rect 4752 6760 4844 6762
rect 4752 6704 4802 6760
rect 4752 6702 4844 6704
rect 4797 6700 4844 6702
rect 4908 6700 4914 6764
rect 5625 6762 5691 6765
rect 11421 6762 11487 6765
rect 18045 6762 18111 6765
rect 5625 6760 8218 6762
rect 5625 6704 5630 6760
rect 5686 6704 8218 6760
rect 5625 6702 8218 6704
rect 4797 6699 4863 6700
rect 5625 6699 5691 6702
rect 8158 6626 8218 6702
rect 11421 6760 18111 6762
rect 11421 6704 11426 6760
rect 11482 6704 18050 6760
rect 18106 6704 18111 6760
rect 11421 6702 18111 6704
rect 11421 6699 11487 6702
rect 18045 6699 18111 6702
rect 12433 6626 12499 6629
rect 8158 6624 12499 6626
rect 8158 6568 12438 6624
rect 12494 6568 12499 6624
rect 8158 6566 12499 6568
rect 12433 6563 12499 6566
rect 16113 6626 16179 6629
rect 17350 6626 17356 6628
rect 16113 6624 17356 6626
rect 16113 6568 16118 6624
rect 16174 6568 17356 6624
rect 16113 6566 17356 6568
rect 16113 6563 16179 6566
rect 17350 6564 17356 6566
rect 17420 6564 17426 6628
rect 18413 6626 18479 6629
rect 19200 6626 20000 6656
rect 18413 6624 20000 6626
rect 18413 6568 18418 6624
rect 18474 6568 20000 6624
rect 18413 6566 20000 6568
rect 18413 6563 18479 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 19200 6536 20000 6566
rect 17606 6495 17922 6496
rect 10501 6490 10567 6493
rect 10685 6490 10751 6493
rect 11697 6490 11763 6493
rect 10501 6488 11763 6490
rect 10501 6432 10506 6488
rect 10562 6432 10690 6488
rect 10746 6432 11702 6488
rect 11758 6432 11763 6488
rect 10501 6430 11763 6432
rect 10501 6427 10567 6430
rect 10685 6427 10751 6430
rect 11697 6427 11763 6430
rect 16614 6428 16620 6492
rect 16684 6490 16690 6492
rect 17309 6490 17375 6493
rect 16684 6488 17375 6490
rect 16684 6432 17314 6488
rect 17370 6432 17375 6488
rect 16684 6430 17375 6432
rect 16684 6428 16690 6430
rect 17309 6427 17375 6430
rect 3141 6354 3207 6357
rect 7649 6354 7715 6357
rect 3141 6352 7715 6354
rect 3141 6296 3146 6352
rect 3202 6296 7654 6352
rect 7710 6296 7715 6352
rect 3141 6294 7715 6296
rect 3141 6291 3207 6294
rect 7649 6291 7715 6294
rect 8518 6292 8524 6356
rect 8588 6354 8594 6356
rect 12709 6354 12775 6357
rect 8588 6352 12775 6354
rect 8588 6296 12714 6352
rect 12770 6296 12775 6352
rect 8588 6294 12775 6296
rect 8588 6292 8594 6294
rect 12709 6291 12775 6294
rect 14181 6354 14247 6357
rect 18229 6354 18295 6357
rect 14181 6352 18295 6354
rect 14181 6296 14186 6352
rect 14242 6296 18234 6352
rect 18290 6296 18295 6352
rect 14181 6294 18295 6296
rect 14181 6291 14247 6294
rect 18229 6291 18295 6294
rect 5349 6218 5415 6221
rect 16849 6218 16915 6221
rect 5349 6216 16915 6218
rect 5349 6160 5354 6216
rect 5410 6160 16854 6216
rect 16910 6160 16915 6216
rect 5349 6158 16915 6160
rect 5349 6155 5415 6158
rect 16849 6155 16915 6158
rect 3734 6020 3740 6084
rect 3804 6082 3810 6084
rect 5349 6082 5415 6085
rect 3804 6080 5415 6082
rect 3804 6024 5354 6080
rect 5410 6024 5415 6080
rect 3804 6022 5415 6024
rect 3804 6020 3810 6022
rect 5349 6019 5415 6022
rect 10225 6082 10291 6085
rect 11094 6082 11100 6084
rect 10225 6080 11100 6082
rect 10225 6024 10230 6080
rect 10286 6024 11100 6080
rect 10225 6022 11100 6024
rect 10225 6019 10291 6022
rect 11094 6020 11100 6022
rect 11164 6082 11170 6084
rect 11164 6022 11714 6082
rect 11164 6020 11170 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 7649 5946 7715 5949
rect 11053 5946 11119 5949
rect 7649 5944 11119 5946
rect 7649 5888 7654 5944
rect 7710 5888 11058 5944
rect 11114 5888 11119 5944
rect 7649 5886 11119 5888
rect 7649 5883 7715 5886
rect 11053 5883 11119 5886
rect 7414 5748 7420 5812
rect 7484 5810 7490 5812
rect 10777 5810 10843 5813
rect 7484 5808 10843 5810
rect 7484 5752 10782 5808
rect 10838 5752 10843 5808
rect 7484 5750 10843 5752
rect 11654 5810 11714 6022
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 12893 5946 12959 5949
rect 12390 5944 12959 5946
rect 12390 5888 12898 5944
rect 12954 5888 12959 5944
rect 12390 5886 12959 5888
rect 12390 5810 12450 5886
rect 12893 5883 12959 5886
rect 11654 5750 12450 5810
rect 12525 5810 12591 5813
rect 12893 5810 12959 5813
rect 12525 5808 12959 5810
rect 12525 5752 12530 5808
rect 12586 5752 12898 5808
rect 12954 5752 12959 5808
rect 12525 5750 12959 5752
rect 7484 5748 7490 5750
rect 10777 5747 10843 5750
rect 12525 5747 12591 5750
rect 12893 5747 12959 5750
rect 5441 5674 5507 5677
rect 10317 5674 10383 5677
rect 5441 5672 10383 5674
rect 5441 5616 5446 5672
rect 5502 5616 10322 5672
rect 10378 5616 10383 5672
rect 5441 5614 10383 5616
rect 5441 5611 5507 5614
rect 10317 5611 10383 5614
rect 10961 5674 11027 5677
rect 18873 5674 18939 5677
rect 10961 5672 18939 5674
rect 10961 5616 10966 5672
rect 11022 5616 18878 5672
rect 18934 5616 18939 5672
rect 10961 5614 18939 5616
rect 10961 5611 11027 5614
rect 18873 5611 18939 5614
rect 9673 5538 9739 5541
rect 10777 5538 10843 5541
rect 9673 5536 10843 5538
rect 9673 5480 9678 5536
rect 9734 5480 10782 5536
rect 10838 5480 10843 5536
rect 9673 5478 10843 5480
rect 9673 5475 9739 5478
rect 10777 5475 10843 5478
rect 18413 5538 18479 5541
rect 19200 5538 20000 5568
rect 18413 5536 20000 5538
rect 18413 5480 18418 5536
rect 18474 5480 20000 5536
rect 18413 5478 20000 5480
rect 18413 5475 18479 5478
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 19200 5448 20000 5478
rect 17606 5407 17922 5408
rect 10726 5340 10732 5404
rect 10796 5402 10802 5404
rect 10869 5402 10935 5405
rect 12382 5402 12388 5404
rect 10796 5400 12388 5402
rect 10796 5344 10874 5400
rect 10930 5344 12388 5400
rect 10796 5342 12388 5344
rect 10796 5340 10802 5342
rect 10869 5339 10935 5342
rect 12382 5340 12388 5342
rect 12452 5340 12458 5404
rect 9673 5266 9739 5269
rect 16113 5266 16179 5269
rect 9673 5264 16179 5266
rect 9673 5208 9678 5264
rect 9734 5208 16118 5264
rect 16174 5208 16179 5264
rect 9673 5206 16179 5208
rect 9673 5203 9739 5206
rect 16113 5203 16179 5206
rect 5390 5130 5396 5132
rect 1718 5070 5396 5130
rect 0 4994 800 5024
rect 1718 4994 1778 5070
rect 5390 5068 5396 5070
rect 5460 5068 5466 5132
rect 6494 5068 6500 5132
rect 6564 5130 6570 5132
rect 16849 5130 16915 5133
rect 6564 5128 16915 5130
rect 6564 5072 16854 5128
rect 16910 5072 16915 5128
rect 6564 5070 16915 5072
rect 6564 5068 6570 5070
rect 16849 5067 16915 5070
rect 0 4934 1778 4994
rect 7465 4994 7531 4997
rect 9489 4994 9555 4997
rect 7465 4992 9555 4994
rect 7465 4936 7470 4992
rect 7526 4936 9494 4992
rect 9550 4936 9555 4992
rect 7465 4934 9555 4936
rect 0 4904 800 4934
rect 7465 4931 7531 4934
rect 9489 4931 9555 4934
rect 12382 4932 12388 4996
rect 12452 4994 12458 4996
rect 16021 4994 16087 4997
rect 12452 4992 16087 4994
rect 12452 4936 16026 4992
rect 16082 4936 16087 4992
rect 12452 4934 16087 4936
rect 12452 4932 12458 4934
rect 16021 4931 16087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 13813 4858 13879 4861
rect 14222 4858 14228 4860
rect 13813 4856 14228 4858
rect 13813 4800 13818 4856
rect 13874 4800 14228 4856
rect 13813 4798 14228 4800
rect 13813 4795 13879 4798
rect 14222 4796 14228 4798
rect 14292 4796 14298 4860
rect 6678 4660 6684 4724
rect 6748 4722 6754 4724
rect 18229 4722 18295 4725
rect 6748 4720 18295 4722
rect 6748 4664 18234 4720
rect 18290 4664 18295 4720
rect 6748 4662 18295 4664
rect 6748 4660 6754 4662
rect 18229 4659 18295 4662
rect 6310 4524 6316 4588
rect 6380 4586 6386 4588
rect 14917 4586 14983 4589
rect 6380 4584 14983 4586
rect 6380 4528 14922 4584
rect 14978 4528 14983 4584
rect 6380 4526 14983 4528
rect 6380 4524 6386 4526
rect 14917 4523 14983 4526
rect 18413 4450 18479 4453
rect 19200 4450 20000 4480
rect 18413 4448 20000 4450
rect 18413 4392 18418 4448
rect 18474 4392 20000 4448
rect 18413 4390 20000 4392
rect 18413 4387 18479 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 19200 4360 20000 4390
rect 17606 4319 17922 4320
rect 8293 4178 8359 4181
rect 9029 4178 9095 4181
rect 8293 4176 9095 4178
rect 8293 4120 8298 4176
rect 8354 4120 9034 4176
rect 9090 4120 9095 4176
rect 8293 4118 9095 4120
rect 8293 4115 8359 4118
rect 9029 4115 9095 4118
rect 9397 4178 9463 4181
rect 9622 4178 9628 4180
rect 9397 4176 9628 4178
rect 9397 4120 9402 4176
rect 9458 4120 9628 4176
rect 9397 4118 9628 4120
rect 9397 4115 9463 4118
rect 9622 4116 9628 4118
rect 9692 4116 9698 4180
rect 12985 4178 13051 4181
rect 13118 4178 13124 4180
rect 12985 4176 13124 4178
rect 12985 4120 12990 4176
rect 13046 4120 13124 4176
rect 12985 4118 13124 4120
rect 12985 4115 13051 4118
rect 13118 4116 13124 4118
rect 13188 4116 13194 4180
rect 1393 4042 1459 4045
rect 9029 4042 9095 4045
rect 1393 4040 9095 4042
rect 1393 3984 1398 4040
rect 1454 3984 9034 4040
rect 9090 3984 9095 4040
rect 1393 3982 9095 3984
rect 1393 3979 1459 3982
rect 9029 3979 9095 3982
rect 10961 4042 11027 4045
rect 15510 4042 15516 4044
rect 10961 4040 15516 4042
rect 10961 3984 10966 4040
rect 11022 3984 15516 4040
rect 10961 3982 15516 3984
rect 10961 3979 11027 3982
rect 15510 3980 15516 3982
rect 15580 3980 15586 4044
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 11697 3772 11763 3773
rect 11646 3708 11652 3772
rect 11716 3770 11763 3772
rect 11716 3768 11808 3770
rect 11758 3712 11808 3768
rect 11716 3710 11808 3712
rect 11716 3708 11763 3710
rect 11697 3707 11763 3708
rect 5349 3634 5415 3637
rect 17861 3634 17927 3637
rect 5349 3632 17927 3634
rect 5349 3576 5354 3632
rect 5410 3576 17866 3632
rect 17922 3576 17927 3632
rect 5349 3574 17927 3576
rect 5349 3571 5415 3574
rect 17861 3571 17927 3574
rect 9305 3498 9371 3501
rect 16246 3498 16252 3500
rect 9305 3496 16252 3498
rect 9305 3440 9310 3496
rect 9366 3440 16252 3496
rect 9305 3438 16252 3440
rect 9305 3435 9371 3438
rect 16246 3436 16252 3438
rect 16316 3436 16322 3500
rect 18413 3362 18479 3365
rect 19200 3362 20000 3392
rect 18413 3360 20000 3362
rect 18413 3304 18418 3360
rect 18474 3304 20000 3360
rect 18413 3302 20000 3304
rect 18413 3299 18479 3302
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 19200 3272 20000 3302
rect 17606 3231 17922 3232
rect 6269 3090 6335 3093
rect 18137 3090 18203 3093
rect 6269 3088 18203 3090
rect 6269 3032 6274 3088
rect 6330 3032 18142 3088
rect 18198 3032 18203 3088
rect 6269 3030 18203 3032
rect 6269 3027 6335 3030
rect 18137 3027 18203 3030
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 3918 2620 3924 2684
rect 3988 2682 3994 2684
rect 5993 2682 6059 2685
rect 3988 2680 6059 2682
rect 3988 2624 5998 2680
rect 6054 2624 6059 2680
rect 3988 2622 6059 2624
rect 3988 2620 3994 2622
rect 5993 2619 6059 2622
rect 9438 2484 9444 2548
rect 9508 2546 9514 2548
rect 14917 2546 14983 2549
rect 9508 2544 14983 2546
rect 9508 2488 14922 2544
rect 14978 2488 14983 2544
rect 9508 2486 14983 2488
rect 9508 2484 9514 2486
rect 14917 2483 14983 2486
rect 18413 2274 18479 2277
rect 19200 2274 20000 2304
rect 18413 2272 20000 2274
rect 18413 2216 18418 2272
rect 18474 2216 20000 2272
rect 18413 2214 20000 2216
rect 18413 2211 18479 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 19200 2184 20000 2214
rect 17606 2143 17922 2144
<< via3 >>
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 11652 17096 11716 17100
rect 11652 17040 11666 17096
rect 11666 17040 11716 17096
rect 11652 17036 11716 17040
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 9444 15948 9508 16012
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 1716 15268 1780 15332
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 10916 15056 10980 15060
rect 10916 15000 10930 15056
rect 10930 15000 10980 15056
rect 10916 14996 10980 15000
rect 13676 14860 13740 14924
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 5580 14452 5644 14516
rect 12388 14512 12452 14516
rect 12388 14456 12438 14512
rect 12438 14456 12452 14512
rect 12388 14452 12452 14456
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 11100 14044 11164 14108
rect 9628 13908 9692 13972
rect 6684 13832 6748 13836
rect 6684 13776 6734 13832
rect 6734 13776 6748 13832
rect 6684 13772 6748 13776
rect 15516 13772 15580 13836
rect 16252 13772 16316 13836
rect 11468 13636 11532 13700
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 13124 13500 13188 13564
rect 10732 13228 10796 13292
rect 6500 13152 6564 13156
rect 6500 13096 6550 13152
rect 6550 13096 6564 13152
rect 6500 13092 6564 13096
rect 14228 13092 14292 13156
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 7420 12956 7484 13020
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 3924 12820 3988 12884
rect 17356 12820 17420 12884
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 7420 12548 7484 12612
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 15148 12548 15212 12612
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 13308 12276 13372 12340
rect 7420 12004 7484 12068
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 9996 11928 10060 11932
rect 9996 11872 10010 11928
rect 10010 11872 10060 11928
rect 9996 11868 10060 11872
rect 13860 11868 13924 11932
rect 16620 11868 16684 11932
rect 3740 11520 3804 11524
rect 3740 11464 3754 11520
rect 3754 11464 3804 11520
rect 3740 11460 3804 11464
rect 8524 11460 8588 11524
rect 10916 11460 10980 11524
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 9996 11324 10060 11388
rect 11652 11384 11716 11388
rect 11652 11328 11702 11384
rect 11702 11328 11716 11384
rect 11652 11324 11716 11328
rect 14044 11324 14108 11388
rect 11652 11052 11716 11116
rect 13676 11052 13740 11116
rect 9628 10916 9692 10980
rect 17356 10976 17420 10980
rect 17356 10920 17406 10976
rect 17406 10920 17420 10976
rect 17356 10916 17420 10920
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 9628 10840 9692 10844
rect 9628 10784 9642 10840
rect 9642 10784 9692 10840
rect 9628 10780 9692 10784
rect 11100 10780 11164 10844
rect 11652 10780 11716 10844
rect 12388 10840 12452 10844
rect 12388 10784 12438 10840
rect 12438 10784 12452 10840
rect 12388 10780 12452 10784
rect 8340 10508 8404 10572
rect 8708 10372 8772 10436
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 8892 10236 8956 10300
rect 5396 9964 5460 10028
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 5580 9692 5644 9756
rect 6684 9692 6748 9756
rect 10548 9692 10612 9756
rect 9812 9420 9876 9484
rect 11284 9420 11348 9484
rect 8156 9284 8220 9348
rect 9076 9284 9140 9348
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 8892 9148 8956 9212
rect 13860 9012 13924 9076
rect 8156 8876 8220 8940
rect 17356 8876 17420 8940
rect 8340 8740 8404 8804
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 8708 8256 8772 8260
rect 8708 8200 8722 8256
rect 8722 8200 8772 8256
rect 8708 8196 8772 8200
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 9076 8060 9140 8124
rect 14044 7924 14108 7988
rect 11468 7788 11532 7852
rect 11100 7652 11164 7716
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 10548 7516 10612 7580
rect 15148 7244 15212 7308
rect 11284 7168 11348 7172
rect 11284 7112 11334 7168
rect 11334 7112 11348 7168
rect 11284 7108 11348 7112
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 11468 6972 11532 7036
rect 13308 6972 13372 7036
rect 9812 6836 9876 6900
rect 4844 6760 4908 6764
rect 4844 6704 4858 6760
rect 4858 6704 4908 6760
rect 4844 6700 4908 6704
rect 17356 6564 17420 6628
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 16620 6428 16684 6492
rect 8524 6292 8588 6356
rect 3740 6020 3804 6084
rect 11100 6020 11164 6084
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 7420 5748 7484 5812
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 10732 5340 10796 5404
rect 12388 5340 12452 5404
rect 5396 5068 5460 5132
rect 6500 5068 6564 5132
rect 12388 4932 12452 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 14228 4796 14292 4860
rect 6684 4660 6748 4724
rect 6316 4524 6380 4588
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 9628 4116 9692 4180
rect 13124 4116 13188 4180
rect 15516 3980 15580 4044
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 11652 3768 11716 3772
rect 11652 3712 11702 3768
rect 11702 3712 11716 3768
rect 11652 3708 11716 3712
rect 16252 3436 16316 3500
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 3924 2620 3988 2684
rect 9444 2484 9508 2548
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
<< metal4 >>
rect 1944 16896 2264 17456
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1715 15332 1781 15333
rect 1715 15268 1716 15332
rect 1780 15268 1781 15332
rect 1715 15267 1781 15268
rect 1718 6578 1778 15267
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 17440 2924 17456
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 6944 16896 7264 17456
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 5579 14516 5645 14517
rect 5579 14452 5580 14516
rect 5644 14452 5645 14516
rect 5579 14451 5645 14452
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 3739 11524 3805 11525
rect 3739 11460 3740 11524
rect 3804 11460 3805 11524
rect 3739 11459 3805 11460
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 3742 6085 3802 11459
rect 3739 6084 3805 6085
rect 3739 6020 3740 6084
rect 3804 6020 3805 6084
rect 3739 6019 3805 6020
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 3926 2685 3986 12819
rect 4846 6765 4906 11782
rect 5395 10028 5461 10029
rect 5395 9964 5396 10028
rect 5460 9964 5461 10028
rect 5395 9963 5461 9964
rect 4843 6764 4909 6765
rect 4843 6700 4844 6764
rect 4908 6700 4909 6764
rect 4843 6699 4909 6700
rect 5398 5133 5458 9963
rect 5582 9757 5642 14451
rect 6683 13836 6749 13837
rect 6683 13772 6684 13836
rect 6748 13772 6749 13836
rect 6683 13771 6749 13772
rect 6499 13156 6565 13157
rect 6499 13092 6500 13156
rect 6564 13092 6565 13156
rect 6499 13091 6565 13092
rect 6502 12450 6562 13091
rect 6318 12390 6562 12450
rect 5579 9756 5645 9757
rect 5579 9692 5580 9756
rect 5644 9692 5645 9756
rect 5579 9691 5645 9692
rect 5395 5132 5461 5133
rect 5395 5068 5396 5132
rect 5460 5068 5461 5132
rect 5395 5067 5461 5068
rect 6318 4589 6378 12390
rect 6686 9890 6746 13771
rect 6502 9830 6746 9890
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 7604 17440 7924 17456
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 11651 17100 11717 17101
rect 11651 17036 11652 17100
rect 11716 17036 11717 17100
rect 11651 17035 11717 17036
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 9443 16012 9509 16013
rect 9443 15948 9444 16012
rect 9508 15948 9509 16012
rect 9443 15947 9509 15948
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7419 13020 7485 13021
rect 7419 12956 7420 13020
rect 7484 12956 7485 13020
rect 7419 12955 7485 12956
rect 7422 12613 7482 12955
rect 7419 12612 7485 12613
rect 7419 12548 7420 12612
rect 7484 12548 7485 12612
rect 7419 12547 7485 12548
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 7419 12068 7485 12069
rect 7419 12004 7420 12068
rect 7484 12004 7485 12068
rect 7419 12003 7485 12004
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6502 5133 6562 9830
rect 6683 9756 6749 9757
rect 6683 9692 6684 9756
rect 6748 9692 6749 9756
rect 6683 9691 6749 9692
rect 6499 5132 6565 5133
rect 6499 5068 6500 5132
rect 6564 5068 6565 5132
rect 6499 5067 6565 5068
rect 6686 4725 6746 9691
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 7422 5813 7482 12003
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 8523 11524 8589 11525
rect 8523 11460 8524 11524
rect 8588 11460 8589 11524
rect 8523 11459 8589 11460
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 8339 10572 8405 10573
rect 8339 10508 8340 10572
rect 8404 10508 8405 10572
rect 8339 10507 8405 10508
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 8155 9348 8221 9349
rect 8155 9284 8156 9348
rect 8220 9284 8221 9348
rect 8155 9283 8221 9284
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 8158 8941 8218 9283
rect 8155 8940 8221 8941
rect 8155 8876 8156 8940
rect 8220 8876 8221 8940
rect 8155 8875 8221 8876
rect 8342 8805 8402 10507
rect 8339 8804 8405 8805
rect 8339 8740 8340 8804
rect 8404 8740 8405 8804
rect 8339 8739 8405 8740
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7419 5812 7485 5813
rect 7419 5748 7420 5812
rect 7484 5748 7485 5812
rect 7419 5747 7485 5748
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6683 4724 6749 4725
rect 6683 4660 6684 4724
rect 6748 4660 6749 4724
rect 6683 4659 6749 4660
rect 6315 4588 6381 4589
rect 6315 4524 6316 4588
rect 6380 4524 6381 4588
rect 6315 4523 6381 4524
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 3923 2684 3989 2685
rect 3923 2620 3924 2684
rect 3988 2620 3989 2684
rect 3923 2619 3989 2620
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 2128 7264 2688
rect 7604 5472 7924 6496
rect 8526 6357 8586 11459
rect 8707 10436 8773 10437
rect 8707 10372 8708 10436
rect 8772 10372 8773 10436
rect 8707 10371 8773 10372
rect 8710 8261 8770 10371
rect 8891 10300 8957 10301
rect 8891 10236 8892 10300
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 8894 9213 8954 10235
rect 9075 9348 9141 9349
rect 9075 9284 9076 9348
rect 9140 9284 9141 9348
rect 9075 9283 9141 9284
rect 8891 9212 8957 9213
rect 8891 9148 8892 9212
rect 8956 9148 8957 9212
rect 8891 9147 8957 9148
rect 8707 8260 8773 8261
rect 8707 8196 8708 8260
rect 8772 8196 8773 8260
rect 8707 8195 8773 8196
rect 9078 8125 9138 9283
rect 9075 8124 9141 8125
rect 9075 8060 9076 8124
rect 9140 8060 9141 8124
rect 9075 8059 9141 8060
rect 8523 6356 8589 6357
rect 8523 6292 8524 6356
rect 8588 6292 8589 6356
rect 8523 6291 8589 6292
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 9446 2549 9506 15947
rect 10915 15060 10981 15061
rect 10915 14996 10916 15060
rect 10980 14996 10981 15060
rect 10915 14995 10981 14996
rect 9627 13972 9693 13973
rect 9627 13908 9628 13972
rect 9692 13908 9693 13972
rect 9627 13907 9693 13908
rect 9630 10981 9690 13907
rect 10731 13292 10797 13293
rect 10731 13228 10732 13292
rect 10796 13228 10797 13292
rect 10731 13227 10797 13228
rect 9995 11932 10061 11933
rect 9995 11868 9996 11932
rect 10060 11868 10061 11932
rect 9995 11867 10061 11868
rect 9998 11389 10058 11867
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 9627 10844 9693 10845
rect 9627 10780 9628 10844
rect 9692 10780 9693 10844
rect 9627 10779 9693 10780
rect 9630 4181 9690 10779
rect 10547 9756 10613 9757
rect 10547 9692 10548 9756
rect 10612 9692 10613 9756
rect 10547 9691 10613 9692
rect 9811 9484 9877 9485
rect 9811 9420 9812 9484
rect 9876 9420 9877 9484
rect 9811 9419 9877 9420
rect 9814 6901 9874 9419
rect 10550 7581 10610 9691
rect 10547 7580 10613 7581
rect 10547 7516 10548 7580
rect 10612 7516 10613 7580
rect 10547 7515 10613 7516
rect 9811 6900 9877 6901
rect 9811 6836 9812 6900
rect 9876 6836 9877 6900
rect 9811 6835 9877 6836
rect 10734 5405 10794 13227
rect 10918 11525 10978 14995
rect 11099 14108 11165 14109
rect 11099 14044 11100 14108
rect 11164 14044 11165 14108
rect 11099 14043 11165 14044
rect 10915 11524 10981 11525
rect 10915 11460 10916 11524
rect 10980 11460 10981 11524
rect 10915 11459 10981 11460
rect 11102 10845 11162 14043
rect 11467 13700 11533 13701
rect 11467 13636 11468 13700
rect 11532 13636 11533 13700
rect 11467 13635 11533 13636
rect 11099 10844 11165 10845
rect 11099 10780 11100 10844
rect 11164 10780 11165 10844
rect 11099 10779 11165 10780
rect 11283 9484 11349 9485
rect 11283 9420 11284 9484
rect 11348 9420 11349 9484
rect 11283 9419 11349 9420
rect 11099 7716 11165 7717
rect 11099 7652 11100 7716
rect 11164 7652 11165 7716
rect 11099 7651 11165 7652
rect 11102 6085 11162 7651
rect 11286 7173 11346 9419
rect 11470 7853 11530 13635
rect 11654 11389 11714 17035
rect 11944 16896 12264 17456
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 12604 17440 12924 17456
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12387 14516 12453 14517
rect 12387 14452 12388 14516
rect 12452 14452 12453 14516
rect 12387 14451 12453 14452
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11651 11388 11717 11389
rect 11651 11324 11652 11388
rect 11716 11324 11717 11388
rect 11651 11323 11717 11324
rect 11654 11117 11714 11323
rect 11651 11116 11717 11117
rect 11651 11052 11652 11116
rect 11716 11052 11717 11116
rect 11651 11051 11717 11052
rect 11651 10844 11717 10845
rect 11651 10780 11652 10844
rect 11716 10780 11717 10844
rect 11651 10779 11717 10780
rect 11467 7852 11533 7853
rect 11467 7788 11468 7852
rect 11532 7788 11533 7852
rect 11467 7787 11533 7788
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 11470 7037 11530 7787
rect 11467 7036 11533 7037
rect 11467 6972 11468 7036
rect 11532 6972 11533 7036
rect 11467 6971 11533 6972
rect 11099 6084 11165 6085
rect 11099 6020 11100 6084
rect 11164 6020 11165 6084
rect 11099 6019 11165 6020
rect 10731 5404 10797 5405
rect 10731 5340 10732 5404
rect 10796 5340 10797 5404
rect 10731 5339 10797 5340
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 11654 3773 11714 10779
rect 11944 10368 12264 11392
rect 12390 10845 12450 14451
rect 12604 14176 12924 15200
rect 16944 16896 17264 17456
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 13675 14924 13741 14925
rect 13675 14860 13676 14924
rect 13740 14860 13741 14924
rect 13675 14859 13741 14860
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 13123 13564 13189 13565
rect 13123 13500 13124 13564
rect 13188 13500 13189 13564
rect 13123 13499 13189 13500
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12387 10844 12453 10845
rect 12387 10780 12388 10844
rect 12452 10780 12453 10844
rect 12387 10779 12453 10780
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12387 5404 12453 5405
rect 12387 5340 12388 5404
rect 12452 5340 12453 5404
rect 12387 5339 12453 5340
rect 12390 4997 12450 5339
rect 12387 4996 12453 4997
rect 12387 4932 12388 4996
rect 12452 4932 12453 4996
rect 12387 4931 12453 4932
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11651 3772 11717 3773
rect 11651 3708 11652 3772
rect 11716 3708 11717 3772
rect 11651 3707 11717 3708
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 9443 2548 9509 2549
rect 9443 2484 9444 2548
rect 9508 2484 9509 2548
rect 9443 2483 9509 2484
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 2128 12264 2688
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 13126 4181 13186 13499
rect 13307 12340 13373 12341
rect 13307 12276 13308 12340
rect 13372 12276 13373 12340
rect 13307 12275 13373 12276
rect 13310 7037 13370 12275
rect 13678 11117 13738 14859
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 15515 13836 15581 13837
rect 15515 13772 15516 13836
rect 15580 13772 15581 13836
rect 15515 13771 15581 13772
rect 16251 13836 16317 13837
rect 16251 13772 16252 13836
rect 16316 13772 16317 13836
rect 16251 13771 16317 13772
rect 14227 13156 14293 13157
rect 14227 13092 14228 13156
rect 14292 13092 14293 13156
rect 14227 13091 14293 13092
rect 13859 11932 13925 11933
rect 13859 11868 13860 11932
rect 13924 11868 13925 11932
rect 13859 11867 13925 11868
rect 13675 11116 13741 11117
rect 13675 11052 13676 11116
rect 13740 11052 13741 11116
rect 13675 11051 13741 11052
rect 13862 9077 13922 11867
rect 14043 11388 14109 11389
rect 14043 11324 14044 11388
rect 14108 11324 14109 11388
rect 14043 11323 14109 11324
rect 13859 9076 13925 9077
rect 13859 9012 13860 9076
rect 13924 9012 13925 9076
rect 13859 9011 13925 9012
rect 14046 7989 14106 11323
rect 14043 7988 14109 7989
rect 14043 7924 14044 7988
rect 14108 7924 14109 7988
rect 14043 7923 14109 7924
rect 13307 7036 13373 7037
rect 13307 6972 13308 7036
rect 13372 6972 13373 7036
rect 13307 6971 13373 6972
rect 14230 4861 14290 13091
rect 15147 12612 15213 12613
rect 15147 12548 15148 12612
rect 15212 12548 15213 12612
rect 15147 12547 15213 12548
rect 15150 7309 15210 12547
rect 15147 7308 15213 7309
rect 15147 7244 15148 7308
rect 15212 7244 15213 7308
rect 15147 7243 15213 7244
rect 14227 4860 14293 4861
rect 14227 4796 14228 4860
rect 14292 4796 14293 4860
rect 14227 4795 14293 4796
rect 13123 4180 13189 4181
rect 13123 4116 13124 4180
rect 13188 4116 13189 4180
rect 13123 4115 13189 4116
rect 15518 4045 15578 13771
rect 15515 4044 15581 4045
rect 15515 3980 15516 4044
rect 15580 3980 15581 4044
rect 15515 3979 15581 3980
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 16254 3501 16314 13771
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 17604 17440 17924 17456
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17355 12884 17421 12885
rect 17355 12820 17356 12884
rect 17420 12820 17421 12884
rect 17355 12819 17421 12820
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 17358 10981 17418 12819
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17355 10980 17421 10981
rect 17355 10916 17356 10980
rect 17420 10916 17421 10980
rect 17355 10915 17421 10916
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17355 8940 17421 8941
rect 17355 8876 17356 8940
rect 17420 8876 17421 8940
rect 17355 8875 17421 8876
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 17358 6629 17418 8875
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17355 6628 17421 6629
rect 17355 6564 17356 6628
rect 17420 6564 17421 6628
rect 17355 6563 17421 6564
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16251 3500 16317 3501
rect 16251 3436 16252 3500
rect 16316 3436 16317 3500
rect 16251 3435 16317 3436
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
<< via4 >>
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1630 6342 1866 6578
rect 1986 3058 2222 3294
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 4758 11782 4994 12018
rect 6986 13058 7222 13294
rect 7646 13718 7882 13954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
rect 11986 13058 12222 13294
rect 12646 13718 12882 13954
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 11986 3058 12222 3294
rect 12646 3718 12882 3954
rect 16986 13058 17222 13294
rect 17646 13718 17882 13954
rect 16534 11932 16770 12018
rect 16534 11868 16620 11932
rect 16620 11868 16684 11932
rect 16684 11868 16770 11932
rect 16534 11782 16770 11868
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16534 6492 16770 6578
rect 16534 6428 16620 6492
rect 16620 6428 16684 6492
rect 16684 6428 16770 6492
rect 16534 6342 16770 6428
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 16986 3058 17222 3294
rect 17646 3718 17882 3954
<< metal5 >>
rect 1056 13954 18908 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 18908 13954
rect 1056 13676 18908 13718
rect 1056 13294 18908 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 18908 13294
rect 1056 13016 18908 13058
rect 4716 12018 16812 12060
rect 4716 11782 4758 12018
rect 4994 11782 16534 12018
rect 16770 11782 16812 12018
rect 4716 11740 16812 11782
rect 1056 8954 18908 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 18908 8954
rect 1056 8676 18908 8718
rect 1056 8294 18908 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 18908 8294
rect 1056 8016 18908 8058
rect 1588 6578 16812 6620
rect 1588 6342 1630 6578
rect 1866 6342 16534 6578
rect 16770 6342 16812 6578
rect 1588 6300 16812 6342
rect 1056 3954 18908 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 18908 3954
rect 1056 3676 18908 3718
rect 1056 3294 18908 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 18908 3294
rect 1056 3016 18908 3058
use sky130_fd_sc_hd__and3_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 1704896540
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _167_
timestamp 1704896540
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1704896540
transform -1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _173_
timestamp 1704896540
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _174_
timestamp 1704896540
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7912 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5152 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _180_
timestamp 1704896540
transform -1 0 12788 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18492 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _183_
timestamp 1704896540
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _185_
timestamp 1704896540
transform -1 0 15640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_2  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1704896540
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 1704896540
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1704896540
transform -1 0 14352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4692 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _193_
timestamp 1704896540
transform -1 0 14260 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1704896540
transform -1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 1704896540
transform -1 0 6072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 1704896540
transform -1 0 11408 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12144 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15272 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1704896540
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _203_
timestamp 1704896540
transform 1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1704896540
transform 1 0 7268 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 1704896540
transform -1 0 8924 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1704896540
transform -1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _207_
timestamp 1704896540
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _208_
timestamp 1704896540
transform -1 0 9752 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _210_
timestamp 1704896540
transform 1 0 10488 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _211_
timestamp 1704896540
transform -1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _212_
timestamp 1704896540
transform -1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1704896540
transform -1 0 4784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1704896540
transform 1 0 5704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1704896540
transform -1 0 12972 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _217_
timestamp 1704896540
transform 1 0 7268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _218_
timestamp 1704896540
transform 1 0 10580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1704896540
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _220_
timestamp 1704896540
transform 1 0 12328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _221_
timestamp 1704896540
transform -1 0 5704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _222_
timestamp 1704896540
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _223_
timestamp 1704896540
transform -1 0 13984 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp 1704896540
transform 1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _225_
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1704896540
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _227_
timestamp 1704896540
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _229_
timestamp 1704896540
transform -1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _230_
timestamp 1704896540
transform -1 0 15364 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 1704896540
transform 1 0 4784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _232_
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1704896540
transform -1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _234_
timestamp 1704896540
transform -1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 1704896540
transform -1 0 18308 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1704896540
transform -1 0 2852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1704896540
transform -1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp 1704896540
transform -1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _241_
timestamp 1704896540
transform -1 0 8096 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _242_
timestamp 1704896540
transform 1 0 3864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1704896540
transform 1 0 11408 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _244_
timestamp 1704896540
transform -1 0 3312 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _245_
timestamp 1704896540
transform -1 0 2576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17204 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _247_
timestamp 1704896540
transform -1 0 14996 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _248_
timestamp 1704896540
transform -1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _249_
timestamp 1704896540
transform 1 0 2208 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1704896540
transform -1 0 6624 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _252_
timestamp 1704896540
transform 1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1704896540
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _254_
timestamp 1704896540
transform 1 0 14904 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _257_
timestamp 1704896540
transform -1 0 4508 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _258_
timestamp 1704896540
transform -1 0 13248 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1704896540
transform -1 0 3588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 1704896540
transform -1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1704896540
transform 1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1704896540
transform -1 0 14628 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1704896540
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _264_
timestamp 1704896540
transform 1 0 2576 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1704896540
transform -1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1704896540
transform -1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _267_
timestamp 1704896540
transform -1 0 14720 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _268_
timestamp 1704896540
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1704896540
transform -1 0 13432 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _270_
timestamp 1704896540
transform -1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _271_
timestamp 1704896540
transform -1 0 11960 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1704896540
transform 1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1704896540
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _274_
timestamp 1704896540
transform -1 0 14720 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11592 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _276_
timestamp 1704896540
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _277_
timestamp 1704896540
transform 1 0 11684 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _278_
timestamp 1704896540
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _279_
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 1704896540
transform 1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _281_
timestamp 1704896540
transform -1 0 17572 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1704896540
transform -1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp 1704896540
transform 1 0 5704 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _284_
timestamp 1704896540
transform -1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _286_
timestamp 1704896540
transform -1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15824 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 1704896540
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _289_
timestamp 1704896540
transform -1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2300 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _291_
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _292_
timestamp 1704896540
transform 1 0 13156 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _293_
timestamp 1704896540
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1704896540
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1704896540
transform -1 0 16192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1704896540
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1704896540
transform 1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1704896540
transform -1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1704896540
transform -1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1704896540
transform -1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1704896540
transform -1 0 15364 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1704896540
transform -1 0 11408 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1704896540
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1704896540
transform -1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1704896540
transform 1 0 14628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1704896540
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1704896540
transform -1 0 17204 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1704896540
transform -1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1704896540
transform -1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1704896540
transform 1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1704896540
transform -1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1704896540
transform 1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1704896540
transform -1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _317_
timestamp 1704896540
transform 1 0 2668 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1704896540
transform 1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1704896540
transform -1 0 11040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1704896540
transform -1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1704896540
transform -1 0 7268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1704896540
transform 1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1704896540
transform -1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1704896540
transform 1 0 13248 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1704896540
transform 1 0 3128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1704896540
transform -1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1704896540
transform 1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _331_
timestamp 1704896540
transform 1 0 11684 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1704896540
transform 1 0 6532 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1704896540
transform -1 0 6532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1704896540
transform 1 0 11960 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1704896540
transform -1 0 13340 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _338_
timestamp 1704896540
transform -1 0 8464 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1704896540
transform 1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _340_
timestamp 1704896540
transform -1 0 9752 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _341_
timestamp 1704896540
transform 1 0 16008 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _342_
timestamp 1704896540
transform -1 0 5980 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _343_
timestamp 1704896540
transform 1 0 3956 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _344_
timestamp 1704896540
transform 1 0 9476 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _345_
timestamp 1704896540
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _346_
timestamp 1704896540
transform 1 0 6716 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _347_
timestamp 1704896540
transform -1 0 6256 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _348_
timestamp 1704896540
transform 1 0 11868 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _349_
timestamp 1704896540
transform 1 0 9568 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _350_
timestamp 1704896540
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp 1704896540
transform -1 0 12604 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp 1704896540
transform 1 0 2668 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _353_
timestamp 1704896540
transform 1 0 8372 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _354_
timestamp 1704896540
transform 1 0 2392 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _355_
timestamp 1704896540
transform 1 0 4784 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 1704896540
transform 1 0 13524 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _357_
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _358_
timestamp 1704896540
transform 1 0 15272 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _359_
timestamp 1704896540
transform 1 0 2944 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _360_
timestamp 1704896540
transform 1 0 8004 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _361_
timestamp 1704896540
transform 1 0 3956 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_1  _370_
timestamp 1704896540
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform -1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1704896540
transform -1 0 2024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1704896540
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1704896540
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1704896540
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 1704896540
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__C
timestamp 1704896540
transform -1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1704896540
transform 1 0 10212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__B
timestamp 1704896540
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1704896540
transform -1 0 3128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__B
timestamp 1704896540
transform -1 0 2944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1704896540
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B
timestamp 1704896540
transform 1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1704896540
transform -1 0 17296 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1704896540
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A1_N
timestamp 1704896540
transform 1 0 10028 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__B1
timestamp 1704896540
transform -1 0 11868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__B2
timestamp 1704896540
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1704896540
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A1
timestamp 1704896540
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A2
timestamp 1704896540
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__B1
timestamp 1704896540
transform 1 0 5428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1704896540
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A1
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__B1
timestamp 1704896540
transform 1 0 10672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A2
timestamp 1704896540
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1704896540
transform 1 0 17572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A1
timestamp 1704896540
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A2
timestamp 1704896540
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__B1
timestamp 1704896540
transform 1 0 8096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B
timestamp 1704896540
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__C
timestamp 1704896540
transform 1 0 12788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__D
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1704896540
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1704896540
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B
timestamp 1704896540
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__C
timestamp 1704896540
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__D
timestamp 1704896540
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1704896540
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__B
timestamp 1704896540
transform -1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A_N
timestamp 1704896540
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__B
timestamp 1704896540
transform 1 0 17940 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__C
timestamp 1704896540
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__D
timestamp 1704896540
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A_N
timestamp 1704896540
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__B
timestamp 1704896540
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__D
timestamp 1704896540
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A1
timestamp 1704896540
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A2
timestamp 1704896540
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__B
timestamp 1704896540
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A1
timestamp 1704896540
transform -1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1704896540
transform 1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B
timestamp 1704896540
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1704896540
transform -1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__B
timestamp 1704896540
transform -1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1704896540
transform 1 0 4876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__B
timestamp 1704896540
transform 1 0 5244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1704896540
transform -1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1704896540
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 1704896540
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__C
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A1
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A2
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__B1
timestamp 1704896540
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B
timestamp 1704896540
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A1
timestamp 1704896540
transform 1 0 12420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A2
timestamp 1704896540
transform 1 0 12972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A3
timestamp 1704896540
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A_N
timestamp 1704896540
transform -1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__B
timestamp 1704896540
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1704896540
transform 1 0 7544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B
timestamp 1704896540
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B
timestamp 1704896540
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1704896540
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A2
timestamp 1704896540
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__C
timestamp 1704896540
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1704896540
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1704896540
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__C1
timestamp 1704896540
transform 1 0 13892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1704896540
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1704896540
transform 1 0 13156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1704896540
transform 1 0 8464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__B
timestamp 1704896540
transform -1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B
timestamp 1704896540
transform -1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1704896540
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A2
timestamp 1704896540
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B
timestamp 1704896540
transform -1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__C
timestamp 1704896540
transform -1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1704896540
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__C
timestamp 1704896540
transform 1 0 16652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1704896540
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B
timestamp 1704896540
transform -1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1704896540
transform -1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B
timestamp 1704896540
transform -1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1704896540
transform -1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1
timestamp 1704896540
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A2
timestamp 1704896540
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B1
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1704896540
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B
timestamp 1704896540
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__C
timestamp 1704896540
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1704896540
transform 1 0 4692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__C
timestamp 1704896540
transform 1 0 4324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1704896540
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B
timestamp 1704896540
transform 1 0 15548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1704896540
transform -1 0 4784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 1704896540
transform -1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1704896540
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1704896540
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1704896540
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A2
timestamp 1704896540
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B1
timestamp 1704896540
transform -1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1704896540
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B
timestamp 1704896540
transform -1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__C
timestamp 1704896540
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1704896540
transform 1 0 17664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__C
timestamp 1704896540
transform -1 0 17664 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1704896540
transform 1 0 3036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1704896540
transform 1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__B
timestamp 1704896540
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1704896540
transform -1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1704896540
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__C
timestamp 1704896540
transform -1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1704896540
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1704896540
transform 1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B
timestamp 1704896540
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__D
timestamp 1704896540
transform -1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A2
timestamp 1704896540
transform -1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B1
timestamp 1704896540
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__C1
timestamp 1704896540
transform -1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1704896540
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B
timestamp 1704896540
transform 1 0 14536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1704896540
transform -1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1704896540
transform 1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1704896540
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1704896540
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1704896540
transform -1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__B
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A1
timestamp 1704896540
transform 1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A2
timestamp 1704896540
transform 1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A3
timestamp 1704896540
transform 1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B1
timestamp 1704896540
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__B1
timestamp 1704896540
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__C1
timestamp 1704896540
transform 1 0 7268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A1
timestamp 1704896540
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A2
timestamp 1704896540
transform 1 0 16100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A3
timestamp 1704896540
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A4
timestamp 1704896540
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B1
timestamp 1704896540
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1704896540
transform 1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__B
timestamp 1704896540
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__C
timestamp 1704896540
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__D
timestamp 1704896540
transform -1 0 3864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1704896540
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B
timestamp 1704896540
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1704896540
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1704896540
transform 1 0 15916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__C
timestamp 1704896540
transform 1 0 14996 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__B
timestamp 1704896540
transform -1 0 14996 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__B
timestamp 1704896540
transform 1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1704896540
transform 1 0 3036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__B
timestamp 1704896540
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__C
timestamp 1704896540
transform -1 0 3588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__C
timestamp 1704896540
transform -1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__D
timestamp 1704896540
transform -1 0 13892 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2
timestamp 1704896540
transform -1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__C1
timestamp 1704896540
transform -1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1704896540
transform -1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1704896540
transform -1 0 16008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1704896540
transform 1 0 12144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B
timestamp 1704896540
transform -1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B2
timestamp 1704896540
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__C1
timestamp 1704896540
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 1704896540
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B
timestamp 1704896540
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1704896540
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1704896540
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1704896540
transform -1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1704896540
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A1
timestamp 1704896540
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A2
timestamp 1704896540
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__B1
timestamp 1704896540
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1704896540
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__B
timestamp 1704896540
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A_N
timestamp 1704896540
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__B
timestamp 1704896540
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__C
timestamp 1704896540
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A1
timestamp 1704896540
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A2
timestamp 1704896540
transform -1 0 15364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__D1
timestamp 1704896540
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__B
timestamp 1704896540
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 1704896540
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A2
timestamp 1704896540
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1704896540
transform 1 0 3404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__B
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__C
timestamp 1704896540
transform 1 0 2300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1704896540
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__B
timestamp 1704896540
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A1
timestamp 1704896540
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A2
timestamp 1704896540
transform -1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1704896540
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1704896540
transform -1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A
timestamp 1704896540
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1704896540
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1704896540
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1704896540
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1704896540
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1704896540
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1704896540
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A
timestamp 1704896540
transform 1 0 18032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 1704896540
transform -1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1704896540
transform 1 0 10488 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1704896540
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1704896540
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1704896540
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1704896540
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1704896540
transform -1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1704896540
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1704896540
transform 1 0 13064 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1704896540
transform 1 0 7636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1704896540
transform 1 0 15456 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1704896540
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1704896540
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 1704896540
transform -1 0 2576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1704896540
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1704896540
transform -1 0 17848 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1704896540
transform -1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 1704896540
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1704896540
transform 1 0 3404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1704896540
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1704896540
transform -1 0 13892 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1704896540
transform 1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1704896540
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1704896540
transform 1 0 15824 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__D
timestamp 1704896540
transform -1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__D
timestamp 1704896540
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__D
timestamp 1704896540
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1704896540
transform -1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1704896540
transform -1 0 8832 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1704896540
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold2_A
timestamp 1704896540
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1704896540
transform -1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output2_A
timestamp 1704896540
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1704896540
transform -1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9200 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 8096 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 12696 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  clkload1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  clkload2
timestamp 1704896540
transform 1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 1704896540
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_61
timestamp 1704896540
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1704896540
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_89
timestamp 1704896540
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_145
timestamp 1704896540
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1704896540
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_185
timestamp 1704896540
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_85
timestamp 1704896540
transform 1 0 8924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_97
timestamp 1704896540
transform 1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_107
timestamp 1704896540
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_121
timestamp 1704896540
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_129
timestamp 1704896540
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_133
timestamp 1704896540
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_145
timestamp 1704896540
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_148
timestamp 1704896540
transform 1 0 14720 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_152
timestamp 1704896540
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_164
timestamp 1704896540
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1704896540
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_11
timestamp 1704896540
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_19
timestamp 1704896540
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1704896540
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_90
timestamp 1704896540
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_123
timestamp 1704896540
transform 1 0 12420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_127
timestamp 1704896540
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_131
timestamp 1704896540
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_184
timestamp 1704896540
transform 1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_19
timestamp 1704896540
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1704896540
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_60
timestamp 1704896540
transform 1 0 6624 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_66
timestamp 1704896540
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_77
timestamp 1704896540
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_85
timestamp 1704896540
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_118
timestamp 1704896540
transform 1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_122
timestamp 1704896540
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_126
timestamp 1704896540
transform 1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_134
timestamp 1704896540
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_138
timestamp 1704896540
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 1704896540
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 1704896540
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_177
timestamp 1704896540
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_180
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_32
timestamp 1704896540
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 1704896540
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 1704896540
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_60
timestamp 1704896540
transform 1 0 6624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_67
timestamp 1704896540
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_71
timestamp 1704896540
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_75
timestamp 1704896540
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_78
timestamp 1704896540
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_106
timestamp 1704896540
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_111
timestamp 1704896540
transform 1 0 11316 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_119
timestamp 1704896540
transform 1 0 12052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_122
timestamp 1704896540
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_129
timestamp 1704896540
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_145
timestamp 1704896540
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_148
timestamp 1704896540
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_155
timestamp 1704896540
transform 1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_159
timestamp 1704896540
transform 1 0 15732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_169
timestamp 1704896540
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_178
timestamp 1704896540
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_182
timestamp 1704896540
transform 1 0 17848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1704896540
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_19
timestamp 1704896540
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_23
timestamp 1704896540
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_35
timestamp 1704896540
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_47
timestamp 1704896540
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_65
timestamp 1704896540
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_74
timestamp 1704896540
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_102
timestamp 1704896540
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_106
timestamp 1704896540
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_133
timestamp 1704896540
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_141
timestamp 1704896540
transform 1 0 14076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_153
timestamp 1704896540
transform 1 0 15180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1704896540
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_177
timestamp 1704896540
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_183
timestamp 1704896540
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_187
timestamp 1704896540
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_19
timestamp 1704896540
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_23
timestamp 1704896540
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_44
timestamp 1704896540
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_48
timestamp 1704896540
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_52
timestamp 1704896540
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_64
timestamp 1704896540
transform 1 0 6992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_72
timestamp 1704896540
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1704896540
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_93
timestamp 1704896540
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_98
timestamp 1704896540
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_102
timestamp 1704896540
transform 1 0 10488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_108
timestamp 1704896540
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_112
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_124
timestamp 1704896540
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_129
timestamp 1704896540
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_141
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_151
timestamp 1704896540
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_155
timestamp 1704896540
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_159
timestamp 1704896540
transform 1 0 15732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_167
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_171
timestamp 1704896540
transform 1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_175
timestamp 1704896540
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_179
timestamp 1704896540
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_183
timestamp 1704896540
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_42
timestamp 1704896540
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_46
timestamp 1704896540
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1704896540
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_97
timestamp 1704896540
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_101
timestamp 1704896540
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_109
timestamp 1704896540
transform 1 0 11132 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_120
timestamp 1704896540
transform 1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_124
timestamp 1704896540
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_128
timestamp 1704896540
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_133
timestamp 1704896540
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1704896540
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_188
timestamp 1704896540
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_23
timestamp 1704896540
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_54
timestamp 1704896540
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_61
timestamp 1704896540
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1704896540
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_81
timestamp 1704896540
transform 1 0 8556 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_95
timestamp 1704896540
transform 1 0 9844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_99
timestamp 1704896540
transform 1 0 10212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_107
timestamp 1704896540
transform 1 0 10948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_132
timestamp 1704896540
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_136
timestamp 1704896540
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1704896540
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_158
timestamp 1704896540
transform 1 0 15640 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_162
timestamp 1704896540
transform 1 0 16008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_170
timestamp 1704896540
transform 1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_175
timestamp 1704896540
transform 1 0 17204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_179
timestamp 1704896540
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_185
timestamp 1704896540
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_11
timestamp 1704896540
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_34
timestamp 1704896540
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_75
timestamp 1704896540
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_79
timestamp 1704896540
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_91
timestamp 1704896540
transform 1 0 9476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_104
timestamp 1704896540
transform 1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_133
timestamp 1704896540
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_141
timestamp 1704896540
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_144
timestamp 1704896540
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_148
timestamp 1704896540
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_152
timestamp 1704896540
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_164
timestamp 1704896540
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_172
timestamp 1704896540
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_176
timestamp 1704896540
transform 1 0 17296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_184
timestamp 1704896540
transform 1 0 18032 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1704896540
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_12
timestamp 1704896540
transform 1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_21
timestamp 1704896540
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_32
timestamp 1704896540
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_36
timestamp 1704896540
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 1704896540
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_66
timestamp 1704896540
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 1704896540
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1704896540
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_102
timestamp 1704896540
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_125
timestamp 1704896540
transform 1 0 12604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_129
timestamp 1704896540
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_136
timestamp 1704896540
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_148
timestamp 1704896540
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_152
timestamp 1704896540
transform 1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_164
timestamp 1704896540
transform 1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_172
timestamp 1704896540
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_177
timestamp 1704896540
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_185
timestamp 1704896540
transform 1 0 18124 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_35
timestamp 1704896540
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_43
timestamp 1704896540
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_77
timestamp 1704896540
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_89
timestamp 1704896540
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_92
timestamp 1704896540
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_100
timestamp 1704896540
transform 1 0 10304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_104
timestamp 1704896540
transform 1 0 10672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_108
timestamp 1704896540
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_117
timestamp 1704896540
transform 1 0 11868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_130
timestamp 1704896540
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_134
timestamp 1704896540
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_138
timestamp 1704896540
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_144
timestamp 1704896540
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_148
timestamp 1704896540
transform 1 0 14720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 1704896540
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_180
timestamp 1704896540
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_24
timestamp 1704896540
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_33
timestamp 1704896540
transform 1 0 4140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_45
timestamp 1704896540
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_58
timestamp 1704896540
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_73
timestamp 1704896540
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_79
timestamp 1704896540
transform 1 0 8372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_111
timestamp 1704896540
transform 1 0 11316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_115
timestamp 1704896540
transform 1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1704896540
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_145
timestamp 1704896540
transform 1 0 14444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_157
timestamp 1704896540
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_169
timestamp 1704896540
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_178
timestamp 1704896540
transform 1 0 17480 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp 1704896540
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1704896540
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_61
timestamp 1704896540
transform 1 0 6716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_94
timestamp 1704896540
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_98
timestamp 1704896540
transform 1 0 10120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1704896540
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_120
timestamp 1704896540
transform 1 0 12144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_126
timestamp 1704896540
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_130
timestamp 1704896540
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_142
timestamp 1704896540
transform 1 0 14168 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 1704896540
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1704896540
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1704896540
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_49
timestamp 1704896540
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_56
timestamp 1704896540
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_60
timestamp 1704896540
transform 1 0 6624 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_72
timestamp 1704896540
transform 1 0 7728 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_108
timestamp 1704896540
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_120
timestamp 1704896540
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1704896540
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_177
timestamp 1704896540
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_185
timestamp 1704896540
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_37
timestamp 1704896540
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 1704896540
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_60
timestamp 1704896540
transform 1 0 6624 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_66
timestamp 1704896540
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_72
timestamp 1704896540
transform 1 0 7728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_76
timestamp 1704896540
transform 1 0 8096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_82
timestamp 1704896540
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_87
timestamp 1704896540
transform 1 0 9108 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_91
timestamp 1704896540
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_103
timestamp 1704896540
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_107
timestamp 1704896540
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_121
timestamp 1704896540
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1704896540
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_153
timestamp 1704896540
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1704896540
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_177
timestamp 1704896540
transform 1 0 17388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_189
timestamp 1704896540
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_37
timestamp 1704896540
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_42
timestamp 1704896540
transform 1 0 4968 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_54
timestamp 1704896540
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_63
timestamp 1704896540
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_67
timestamp 1704896540
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_79
timestamp 1704896540
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_92
timestamp 1704896540
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1704896540
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_108
timestamp 1704896540
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_112
timestamp 1704896540
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_116
timestamp 1704896540
transform 1 0 11776 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_147
timestamp 1704896540
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_151
timestamp 1704896540
transform 1 0 14996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_162
timestamp 1704896540
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_166
timestamp 1704896540
transform 1 0 16376 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_179
timestamp 1704896540
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_15
timestamp 1704896540
transform 1 0 2484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_19
timestamp 1704896540
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_23
timestamp 1704896540
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_35
timestamp 1704896540
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_40
timestamp 1704896540
transform 1 0 4784 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1704896540
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_102
timestamp 1704896540
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_106
timestamp 1704896540
transform 1 0 10856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_124
timestamp 1704896540
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_146
timestamp 1704896540
transform 1 0 14536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_154
timestamp 1704896540
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_164
timestamp 1704896540
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1704896540
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1704896540
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_10
timestamp 1704896540
transform 1 0 2024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_17
timestamp 1704896540
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1704896540
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_33
timestamp 1704896540
transform 1 0 4140 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1704896540
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_52
timestamp 1704896540
transform 1 0 5888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1704896540
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_107
timestamp 1704896540
transform 1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_115
timestamp 1704896540
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_119
timestamp 1704896540
transform 1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_123
timestamp 1704896540
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_132
timestamp 1704896540
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_136
timestamp 1704896540
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_150
timestamp 1704896540
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_154
timestamp 1704896540
transform 1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_165
timestamp 1704896540
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_169
timestamp 1704896540
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_178
timestamp 1704896540
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_182
timestamp 1704896540
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_186
timestamp 1704896540
transform 1 0 18216 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_22
timestamp 1704896540
transform 1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_30
timestamp 1704896540
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_42
timestamp 1704896540
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1704896540
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_63
timestamp 1704896540
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_68
timestamp 1704896540
transform 1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_72
timestamp 1704896540
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_105
timestamp 1704896540
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_117
timestamp 1704896540
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_123
timestamp 1704896540
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_135
timestamp 1704896540
transform 1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_140
timestamp 1704896540
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_152
timestamp 1704896540
transform 1 0 15088 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_33
timestamp 1704896540
transform 1 0 4140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_59
timestamp 1704896540
transform 1 0 6532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_64
timestamp 1704896540
transform 1 0 6992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_70
timestamp 1704896540
transform 1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_74
timestamp 1704896540
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_78
timestamp 1704896540
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_104
timestamp 1704896540
transform 1 0 10672 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_116
timestamp 1704896540
transform 1 0 11776 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_128
timestamp 1704896540
transform 1 0 12880 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_132
timestamp 1704896540
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_136
timestamp 1704896540
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_177
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_181
timestamp 1704896540
transform 1 0 17756 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_185
timestamp 1704896540
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_17
timestamp 1704896540
transform 1 0 2668 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_23
timestamp 1704896540
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1704896540
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1704896540
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_73
timestamp 1704896540
transform 1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_77
timestamp 1704896540
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_100
timestamp 1704896540
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_104
timestamp 1704896540
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_118
timestamp 1704896540
transform 1 0 11960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_122
timestamp 1704896540
transform 1 0 12328 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_135
timestamp 1704896540
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1704896540
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_175
timestamp 1704896540
transform 1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_179
timestamp 1704896540
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1704896540
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 1704896540
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_13
timestamp 1704896540
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_23
timestamp 1704896540
transform 1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_34
timestamp 1704896540
transform 1 0 4232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_38
timestamp 1704896540
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_42
timestamp 1704896540
transform 1 0 4968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_50
timestamp 1704896540
transform 1 0 5704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_55
timestamp 1704896540
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1704896540
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1704896540
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_96
timestamp 1704896540
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_108
timestamp 1704896540
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_120
timestamp 1704896540
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_127
timestamp 1704896540
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1704896540
transform 1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_158
timestamp 1704896540
transform 1 0 15640 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_183
timestamp 1704896540
transform 1 0 17940 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_7
timestamp 1704896540
transform 1 0 1748 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_45
timestamp 1704896540
transform 1 0 5244 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1704896540
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_61
timestamp 1704896540
transform 1 0 6716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_73
timestamp 1704896540
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_85
timestamp 1704896540
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_94
timestamp 1704896540
transform 1 0 9752 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_99
timestamp 1704896540
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_117
timestamp 1704896540
transform 1 0 11868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_129
timestamp 1704896540
transform 1 0 12972 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_135
timestamp 1704896540
transform 1 0 13524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_143
timestamp 1704896540
transform 1 0 14260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_148
timestamp 1704896540
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 1704896540
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1704896540
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_33
timestamp 1704896540
transform 1 0 4140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_57
timestamp 1704896540
transform 1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_61
timestamp 1704896540
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_67
timestamp 1704896540
transform 1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 1704896540
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_99
timestamp 1704896540
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_106
timestamp 1704896540
transform 1 0 10856 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_118
timestamp 1704896540
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_122
timestamp 1704896540
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_134
timestamp 1704896540
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_148
timestamp 1704896540
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_152
timestamp 1704896540
transform 1 0 15088 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_155
timestamp 1704896540
transform 1 0 15364 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_167
timestamp 1704896540
transform 1 0 16468 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_179
timestamp 1704896540
transform 1 0 17572 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_15
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_19
timestamp 1704896540
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_22
timestamp 1704896540
transform 1 0 3128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_30
timestamp 1704896540
transform 1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_133
timestamp 1704896540
transform 1 0 13340 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_141
timestamp 1704896540
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_147
timestamp 1704896540
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1704896540
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_189
timestamp 1704896540
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_18
timestamp 1704896540
transform 1 0 2760 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 1704896540
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1704896540
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_43
timestamp 1704896540
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_47
timestamp 1704896540
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_54
timestamp 1704896540
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_58
timestamp 1704896540
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_67
timestamp 1704896540
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1704896540
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_109
timestamp 1704896540
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_125
timestamp 1704896540
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_129
timestamp 1704896540
transform 1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_135
timestamp 1704896540
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1704896540
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_147
timestamp 1704896540
transform 1 0 14628 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_151
timestamp 1704896540
transform 1 0 14996 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_155
timestamp 1704896540
transform 1 0 15364 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_167
timestamp 1704896540
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_179
timestamp 1704896540
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_20
timestamp 1704896540
transform 1 0 2944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_29
timestamp 1704896540
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_33
timestamp 1704896540
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_43
timestamp 1704896540
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1704896540
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_65
timestamp 1704896540
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_77
timestamp 1704896540
transform 1 0 8188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1704896540
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1704896540
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1704896540
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_138
timestamp 1704896540
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_141
timestamp 1704896540
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_149
timestamp 1704896540
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_153
timestamp 1704896540
transform 1 0 15180 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_159
timestamp 1704896540
transform 1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1704896540
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6808 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 9752 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1704896540
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1704896540
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1704896540
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1704896540
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1704896540
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1704896540
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1704896540
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 1704896540
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1704896540
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1704896540
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_10
timestamp 1704896540
transform -1 0 18584 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_11
timestamp 1704896540
transform -1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_12
timestamp 1704896540
transform -1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_13
timestamp 1704896540
transform -1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_14
timestamp 1704896540
transform -1 0 18584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_15
timestamp 1704896540
transform -1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_16
timestamp 1704896540
transform -1 0 18584 0 1 10880
box -38 -48 314 592
<< labels >>
flabel metal4 s 2604 2128 2924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3676 18908 3996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8676 18908 8996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13676 18908 13996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11944 2128 12264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16944 2128 17264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 18908 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 18908 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 13016 18908 13336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 19200 17416 20000 17536 0 FreeSans 480 0 0 0 an[0]
port 2 nsew signal output
flabel metal3 s 19200 16328 20000 16448 0 FreeSans 480 0 0 0 an[1]
port 3 nsew signal output
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 an[2]
port 4 nsew signal output
flabel metal3 s 19200 14152 20000 14272 0 FreeSans 480 0 0 0 an[3]
port 5 nsew signal output
flabel metal3 s 19200 13064 20000 13184 0 FreeSans 480 0 0 0 an[4]
port 6 nsew signal output
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 an[5]
port 7 nsew signal output
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 480 0 0 0 an[6]
port 8 nsew signal output
flabel metal3 s 19200 9800 20000 9920 0 FreeSans 480 0 0 0 an[7]
port 9 nsew signal output
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 clk
port 10 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 rst
port 11 nsew signal input
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 seg[0]
port 12 nsew signal output
flabel metal3 s 19200 7624 20000 7744 0 FreeSans 480 0 0 0 seg[1]
port 13 nsew signal output
flabel metal3 s 19200 6536 20000 6656 0 FreeSans 480 0 0 0 seg[2]
port 14 nsew signal output
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 seg[3]
port 15 nsew signal output
flabel metal3 s 19200 4360 20000 4480 0 FreeSans 480 0 0 0 seg[4]
port 16 nsew signal output
flabel metal3 s 19200 3272 20000 3392 0 FreeSans 480 0 0 0 seg[5]
port 17 nsew signal output
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 seg[6]
port 18 nsew signal output
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel metal1 9982 16864 9982 16864 0 VPWR
rlabel metal1 6808 13158 6808 13158 0 _000_
rlabel metal2 15962 13991 15962 13991 0 _001_
rlabel metal1 6854 12172 6854 12172 0 _002_
rlabel metal1 17802 4794 17802 4794 0 _003_
rlabel metal1 4140 6698 4140 6698 0 _004_
rlabel metal1 9476 2346 9476 2346 0 _005_
rlabel metal2 2162 15351 2162 15351 0 _006_
rlabel metal1 6164 3434 6164 3434 0 _007_
rlabel metal1 10534 10574 10534 10574 0 _008_
rlabel metal2 10902 16031 10902 16031 0 _009_
rlabel metal2 9890 7548 9890 7548 0 _010_
rlabel metal1 5658 13158 5658 13158 0 _011_
rlabel metal3 14191 13124 14191 13124 0 _012_
rlabel metal2 12650 8364 12650 8364 0 _013_
rlabel metal1 7360 6630 7360 6630 0 _014_
rlabel metal1 8740 11662 8740 11662 0 _015_
rlabel metal2 2622 10608 2622 10608 0 _016_
rlabel metal2 5106 9520 5106 9520 0 _017_
rlabel metal2 7866 8075 7866 8075 0 _018_
rlabel metal2 16238 12665 16238 12665 0 _019_
rlabel metal1 2024 7514 2024 7514 0 _020_
rlabel metal1 6808 11322 6808 11322 0 _021_
rlabel metal1 8648 10778 8648 10778 0 _022_
rlabel metal1 8510 11560 8510 11560 0 _023_
rlabel metal1 14582 11016 14582 11016 0 _024_
rlabel metal2 17342 14433 17342 14433 0 _025_
rlabel via2 16882 6171 16882 6171 0 _026_
rlabel via2 1978 8381 1978 8381 0 _027_
rlabel metal2 1794 3536 1794 3536 0 _028_
rlabel metal1 16054 11764 16054 11764 0 _029_
rlabel metal2 18078 9775 18078 9775 0 _030_
rlabel metal1 2162 5338 2162 5338 0 _031_
rlabel metal1 7682 7514 7682 7514 0 _032_
rlabel metal2 5198 13532 5198 13532 0 _033_
rlabel metal1 15417 8874 15417 8874 0 _034_
rlabel metal2 15226 15640 15226 15640 0 _035_
rlabel metal1 7873 14314 7873 14314 0 _036_
rlabel metal2 18170 3485 18170 3485 0 _037_
rlabel metal1 9568 13838 9568 13838 0 _038_
rlabel metal1 15824 12410 15824 12410 0 _039_
rlabel metal2 14674 16830 14674 16830 0 _040_
rlabel metal3 16859 11900 16859 11900 0 _041_
rlabel metal1 12105 2346 12105 2346 0 _042_
rlabel metal1 3871 15470 3871 15470 0 _043_
rlabel metal2 17434 4335 17434 4335 0 _044_
rlabel metal2 12006 14246 12006 14246 0 _045_
rlabel metal1 7406 13838 7406 13838 0 _046_
rlabel metal3 15663 13804 15663 13804 0 _047_
rlabel metal1 13110 15504 13110 15504 0 _048_
rlabel metal1 7544 8058 7544 8058 0 _049_
rlabel metal2 7222 10914 7222 10914 0 _050_
rlabel metal1 10265 11798 10265 11798 0 _051_
rlabel via2 3197 15164 3197 15164 0 _052_
rlabel metal1 4416 3706 4416 3706 0 _053_
rlabel metal4 13340 9656 13340 9656 0 _054_
rlabel metal1 3365 8534 3365 8534 0 _055_
rlabel metal2 13386 16014 13386 16014 0 _056_
rlabel metal1 3772 16422 3772 16422 0 _057_
rlabel metal1 9798 13226 9798 13226 0 _058_
rlabel metal2 16146 5661 16146 5661 0 _059_
rlabel metal2 10258 10727 10258 10727 0 _060_
rlabel metal1 3036 5882 3036 5882 0 _061_
rlabel metal1 7406 3978 7406 3978 0 _062_
rlabel metal1 2208 16762 2208 16762 0 _063_
rlabel metal2 3174 6035 3174 6035 0 _064_
rlabel metal1 2254 16660 2254 16660 0 _065_
rlabel metal1 14582 12716 14582 12716 0 _066_
rlabel metal1 16652 7174 16652 7174 0 _067_
rlabel metal1 13110 13328 13110 13328 0 _068_
rlabel metal1 2530 6970 2530 6970 0 _069_
rlabel metal2 6394 4182 6394 4182 0 _070_
rlabel metal1 4922 14858 4922 14858 0 _071_
rlabel metal2 10166 6460 10166 6460 0 _072_
rlabel metal1 17066 3366 17066 3366 0 _073_
rlabel metal2 9982 4794 9982 4794 0 _074_
rlabel metal1 2576 3910 2576 3910 0 _075_
rlabel metal1 4968 15470 4968 15470 0 _076_
rlabel metal1 13064 4590 13064 4590 0 _077_
rlabel metal2 8142 8228 8142 8228 0 _078_
rlabel metal1 7268 4794 7268 4794 0 _079_
rlabel metal1 10074 9044 10074 9044 0 _080_
rlabel via1 7317 9146 7317 9146 0 _081_
rlabel metal1 10258 4624 10258 4624 0 _082_
rlabel metal2 15042 5610 15042 5610 0 _083_
rlabel metal2 10534 7684 10534 7684 0 _084_
rlabel metal1 2208 7786 2208 7786 0 _085_
rlabel metal3 13041 8364 13041 8364 0 _086_
rlabel metal2 14214 11832 14214 11832 0 _087_
rlabel metal2 14030 15946 14030 15946 0 _088_
rlabel metal2 13938 14093 13938 14093 0 _089_
rlabel metal1 10626 11322 10626 11322 0 _090_
rlabel via2 6026 2635 6026 2635 0 _091_
rlabel metal1 9706 12648 9706 12648 0 _092_
rlabel metal2 17342 4794 17342 4794 0 _093_
rlabel metal4 13892 10472 13892 10472 0 _094_
rlabel metal1 17986 4522 17986 4522 0 _095_
rlabel metal1 8418 3910 8418 3910 0 _096_
rlabel via3 8717 8228 8717 8228 0 _097_
rlabel metal1 6716 11118 6716 11118 0 _098_
rlabel metal1 10028 10506 10028 10506 0 _099_
rlabel metal1 9246 14790 9246 14790 0 _100_
rlabel metal1 13294 5848 13294 5848 0 _101_
rlabel metal1 13846 11118 13846 11118 0 _102_
rlabel metal2 13110 6018 13110 6018 0 _103_
rlabel metal2 9614 15504 9614 15504 0 _104_
rlabel metal2 10626 5202 10626 5202 0 _105_
rlabel metal3 9131 5780 9131 5780 0 _106_
rlabel metal1 18722 14382 18722 14382 0 _107_
rlabel metal2 16974 6595 16974 6595 0 _108_
rlabel metal1 5198 15334 5198 15334 0 _109_
rlabel metal2 12466 3145 12466 3145 0 _110_
rlabel metal3 1955 13396 1955 13396 0 _111_
rlabel metal3 16215 13804 16215 13804 0 _112_
rlabel metal1 3956 12206 3956 12206 0 _113_
rlabel metal1 4830 16524 4830 16524 0 _114_
rlabel via2 14950 4539 14950 4539 0 _115_
rlabel metal1 5804 14042 5804 14042 0 _116_
rlabel metal1 16974 4794 16974 4794 0 _117_
rlabel metal1 18078 3944 18078 3944 0 _118_
rlabel metal2 12834 13464 12834 13464 0 _119_
rlabel metal2 17894 3757 17894 3757 0 _120_
rlabel metal2 4738 13787 4738 13787 0 _121_
rlabel metal1 9506 15538 9506 15538 0 _122_
rlabel metal2 16698 14144 16698 14144 0 _123_
rlabel metal2 3910 14450 3910 14450 0 _124_
rlabel metal2 12650 15742 12650 15742 0 _125_
rlabel metal1 2576 8874 2576 8874 0 _126_
rlabel metal1 6992 7718 6992 7718 0 _127_
rlabel metal1 2346 12410 2346 12410 0 _128_
rlabel metal1 12236 11866 12236 11866 0 _129_
rlabel metal2 4462 11764 4462 11764 0 _130_
rlabel metal2 9522 10948 9522 10948 0 _131_
rlabel metal2 10626 16252 10626 16252 0 _132_
rlabel via2 14950 2533 14950 2533 0 _133_
rlabel metal1 16146 16966 16146 16966 0 _134_
rlabel metal1 14076 15402 14076 15402 0 _135_
rlabel metal1 16376 8058 16376 8058 0 _136_
rlabel metal1 3910 17034 3910 17034 0 _137_
rlabel metal1 12926 17306 12926 17306 0 _138_
rlabel via2 14214 16643 14214 16643 0 _139_
rlabel metal2 13754 7871 13754 7871 0 _140_
rlabel metal1 12190 3536 12190 3536 0 _141_
rlabel metal1 7590 11322 7590 11322 0 _142_
rlabel metal2 13708 7718 13708 7718 0 _143_
rlabel metal2 12742 13651 12742 13651 0 _144_
rlabel metal1 11868 6630 11868 6630 0 _145_
rlabel metal2 8694 13056 8694 13056 0 _146_
rlabel metal1 12006 6800 12006 6800 0 _147_
rlabel metal1 7130 7820 7130 7820 0 _148_
rlabel metal4 14076 9656 14076 9656 0 _149_
rlabel metal1 5934 9962 5934 9962 0 _150_
rlabel metal2 17066 10880 17066 10880 0 _151_
rlabel metal1 17380 11050 17380 11050 0 _152_
rlabel via2 15226 11237 15226 11237 0 _153_
rlabel metal3 4646 8228 4646 8228 0 _154_
rlabel metal1 15870 15028 15870 15028 0 _155_
rlabel metal1 13202 7922 13202 7922 0 _156_
rlabel metal2 2346 12512 2346 12512 0 _157_
rlabel metal1 13662 8058 13662 8058 0 _158_
rlabel metal1 1886 4148 1886 4148 0 _159_
rlabel metal2 13018 7446 13018 7446 0 _160_
rlabel metal1 7222 16592 7222 16592 0 _161_
rlabel metal3 1211 4964 1211 4964 0 clk
rlabel metal1 7498 12138 7498 12138 0 clknet_0_clk
rlabel metal2 8050 4386 8050 4386 0 clknet_2_0__leaf_clk
rlabel metal1 2622 10642 2622 10642 0 clknet_2_1__leaf_clk
rlabel metal1 9338 3978 9338 3978 0 clknet_2_2__leaf_clk
rlabel metal2 13294 16524 13294 16524 0 clknet_2_3__leaf_clk
rlabel metal1 5934 14960 5934 14960 0 decoder.digit\[0\]
rlabel metal1 5658 14790 5658 14790 0 decoder.digit\[1\]
rlabel via2 5474 5661 5474 5661 0 decoder.digit\[2\]
rlabel metal1 2346 16593 2346 16593 0 decoder.digit\[3\]
rlabel metal2 2622 13549 2622 13549 0 net1
rlabel metal2 18538 17391 18538 17391 0 net10
rlabel via2 18538 16405 18538 16405 0 net11
rlabel via2 18538 15317 18538 15317 0 net12
rlabel via2 18262 14229 18262 14229 0 net13
rlabel via2 18538 13141 18538 13141 0 net14
rlabel via2 18538 12053 18538 12053 0 net15
rlabel metal2 18538 10999 18538 10999 0 net16
rlabel metal1 9890 8534 9890 8534 0 net17
rlabel metal1 9108 9078 9108 9078 0 net18
rlabel metal1 16008 9146 16008 9146 0 net2
rlabel metal1 18216 7854 18216 7854 0 net3
rlabel metal1 17940 12410 17940 12410 0 net4
rlabel metal1 16468 12886 16468 12886 0 net5
rlabel metal2 18262 4641 18262 4641 0 net6
rlabel metal3 16376 12716 16376 12716 0 net7
rlabel metal1 18446 2414 18446 2414 0 net8
rlabel metal2 18538 9945 18538 9945 0 net9
rlabel metal1 4646 17272 4646 17272 0 one_second_counter\[0\]
rlabel metal1 8648 6970 8648 6970 0 one_second_counter\[10\]
rlabel metal2 16376 12716 16376 12716 0 one_second_counter\[11\]
rlabel metal1 5520 14382 5520 14382 0 one_second_counter\[12\]
rlabel metal1 18124 13498 18124 13498 0 one_second_counter\[13\]
rlabel metal2 17986 13991 17986 13991 0 one_second_counter\[14\]
rlabel metal1 5014 15674 5014 15674 0 one_second_counter\[15\]
rlabel metal1 9154 3502 9154 3502 0 one_second_counter\[16\]
rlabel metal1 14996 2618 14996 2618 0 one_second_counter\[17\]
rlabel metal1 14904 2482 14904 2482 0 one_second_counter\[18\]
rlabel metal1 17480 13838 17480 13838 0 one_second_counter\[19\]
rlabel metal1 6348 2278 6348 2278 0 one_second_counter\[1\]
rlabel metal1 15640 13838 15640 13838 0 one_second_counter\[20\]
rlabel metal2 15088 13260 15088 13260 0 one_second_counter\[21\]
rlabel metal2 4462 10336 4462 10336 0 one_second_counter\[22\]
rlabel metal1 15180 6834 15180 6834 0 one_second_counter\[23\]
rlabel metal2 6854 7650 6854 7650 0 one_second_counter\[24\]
rlabel metal1 17020 3706 17020 3706 0 one_second_counter\[25\]
rlabel metal1 15272 6426 15272 6426 0 one_second_counter\[26\]
rlabel metal1 5980 2414 5980 2414 0 one_second_counter\[2\]
rlabel metal1 11408 3502 11408 3502 0 one_second_counter\[3\]
rlabel metal2 4738 7344 4738 7344 0 one_second_counter\[4\]
rlabel metal1 9936 15062 9936 15062 0 one_second_counter\[5\]
rlabel metal1 6946 6834 6946 6834 0 one_second_counter\[6\]
rlabel metal1 5290 5814 5290 5814 0 one_second_counter\[7\]
rlabel metal1 12581 4590 12581 4590 0 one_second_counter\[8\]
rlabel metal1 5888 14518 5888 14518 0 one_second_counter\[9\]
rlabel metal1 5980 15062 5980 15062 0 one_second_enable
rlabel via2 1610 15045 1610 15045 0 rst
rlabel via2 18446 8789 18446 8789 0 seg[0]
rlabel via2 18446 7701 18446 7701 0 seg[1]
rlabel via2 18446 6613 18446 6613 0 seg[2]
rlabel via2 18446 5525 18446 5525 0 seg[3]
rlabel via2 18446 4437 18446 4437 0 seg[4]
rlabel via2 18446 3349 18446 3349 0 seg[5]
rlabel via2 18446 2261 18446 2261 0 seg[6]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
